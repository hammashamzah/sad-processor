module template_image_rom(
	input [11:0] addr,
	input clk,
	output out
);
	reg q;

	always @(posedge clk)
	begin
		case(addr)
			12'd00: q <= 1'b1;
			12'd01: q <= 1'b1;
			12'd02: q <= 1'b1;
			12'd03: q <= 1'b1;
			12'd04: q <= 1'b1;
			12'd05: q <= 1'b1;
			12'd06: q <= 1'b1;
			12'd07: q <= 1'b1;
			12'd08: q <= 1'b1;
			12'd09: q <= 1'b1;
			12'd10: q <= 1'b1;
			12'd11: q <= 1'b1;
			12'd12: q <= 1'b1;
			12'd13: q <= 1'b1;
			12'd14: q <= 1'b1;
			12'd15: q <= 1'b1;
			12'd16: q <= 1'b1;
			12'd17: q <= 1'b1;
			12'd18: q <= 1'b1;
			12'd19: q <= 1'b1;
			12'd20: q <= 1'b1;
			12'd21: q <= 1'b1;
			12'd22: q <= 1'b1;
			12'd23: q <= 1'b1;
			12'd24: q <= 1'b1;
			12'd25: q <= 1'b1;
			12'd26: q <= 1'b1;
			12'd27: q <= 1'b1;
			12'd28: q <= 1'b1;
			12'd29: q <= 1'b1;
			12'd30: q <= 1'b1;
			12'd31: q <= 1'b1;
			12'd32: q <= 1'b1;
			12'd33: q <= 1'b1;
			12'd34: q <= 1'b1;
			12'd35: q <= 1'b1;
			12'd36: q <= 1'b1;
			12'd37: q <= 1'b1;
			12'd38: q <= 1'b1;
			12'd39: q <= 1'b1;
			12'd40: q <= 1'b1;
			12'd41: q <= 1'b1;
			12'd42: q <= 1'b1;
			12'd43: q <= 1'b1;
			12'd44: q <= 1'b1;
			12'd45: q <= 1'b1;
			12'd46: q <= 1'b1;
			12'd47: q <= 1'b1;
			12'd48: q <= 1'b1;
			12'd49: q <= 1'b1;
			12'd50: q <= 1'b1;
			12'd51: q <= 1'b1;
			12'd52: q <= 1'b1;
			12'd53: q <= 1'b1;
			12'd54: q <= 1'b1;
			12'd55: q <= 1'b1;
			12'd56: q <= 1'b1;
			12'd57: q <= 1'b1;
			12'd58: q <= 1'b1;
			12'd59: q <= 1'b1;
			12'd60: q <= 1'b1;
			12'd61: q <= 1'b1;
			12'd62: q <= 1'b1;
			12'd63: q <= 1'b1;
			12'd64: q <= 1'b1;
			12'd65: q <= 1'b1;
			12'd66: q <= 1'b1;
			12'd67: q <= 1'b1;
			12'd68: q <= 1'b1;
			12'd69: q <= 1'b1;
			12'd70: q <= 1'b1;
			12'd71: q <= 1'b1;
			12'd72: q <= 1'b1;
			12'd73: q <= 1'b1;
			12'd74: q <= 1'b1;
			12'd75: q <= 1'b1;
			12'd76: q <= 1'b1;
			12'd77: q <= 1'b1;
			12'd78: q <= 1'b1;
			12'd79: q <= 1'b1;
			12'd80: q <= 1'b1;
			12'd81: q <= 1'b1;
			12'd82: q <= 1'b1;
			12'd83: q <= 1'b1;
			12'd84: q <= 1'b1;
			12'd85: q <= 1'b1;
			12'd86: q <= 1'b1;
			12'd87: q <= 1'b1;
			12'd88: q <= 1'b1;
			12'd89: q <= 1'b1;
			12'd90: q <= 1'b1;
			12'd91: q <= 1'b1;
			12'd92: q <= 1'b1;
			12'd93: q <= 1'b1;
			12'd94: q <= 1'b1;
			12'd95: q <= 1'b1;
			12'd96: q <= 1'b1;
			12'd97: q <= 1'b1;
			12'd98: q <= 1'b1;
			12'd99: q <= 1'b1;
			12'd100: q <= 1'b1;
			12'd101: q <= 1'b1;
			12'd102: q <= 1'b1;
			12'd103: q <= 1'b1;
			12'd104: q <= 1'b1;
			12'd105: q <= 1'b1;
			12'd106: q <= 1'b1;
			12'd107: q <= 1'b1;
			12'd108: q <= 1'b1;
			12'd109: q <= 1'b1;
			12'd110: q <= 1'b1;
			12'd111: q <= 1'b1;
			12'd112: q <= 1'b1;
			12'd113: q <= 1'b1;
			12'd114: q <= 1'b1;
			12'd115: q <= 1'b1;
			12'd116: q <= 1'b1;
			12'd117: q <= 1'b1;
			12'd118: q <= 1'b1;
			12'd119: q <= 1'b1;
			12'd120: q <= 1'b1;
			12'd121: q <= 1'b1;
			12'd122: q <= 1'b1;
			12'd123: q <= 1'b1;
			12'd124: q <= 1'b1;
			12'd125: q <= 1'b1;
			12'd126: q <= 1'b1;
			12'd127: q <= 1'b1;
			12'd128: q <= 1'b1;
			12'd129: q <= 1'b1;
			12'd130: q <= 1'b1;
			12'd131: q <= 1'b1;
			12'd132: q <= 1'b1;
			12'd133: q <= 1'b1;
			12'd134: q <= 1'b1;
			12'd135: q <= 1'b1;
			12'd136: q <= 1'b1;
			12'd137: q <= 1'b1;
			12'd138: q <= 1'b1;
			12'd139: q <= 1'b1;
			12'd140: q <= 1'b1;
			12'd141: q <= 1'b1;
			12'd142: q <= 1'b1;
			12'd143: q <= 1'b1;
			12'd144: q <= 1'b1;
			12'd145: q <= 1'b1;
			12'd146: q <= 1'b1;
			12'd147: q <= 1'b1;
			12'd148: q <= 1'b1;
			12'd149: q <= 1'b1;
			12'd150: q <= 1'b1;
			12'd151: q <= 1'b1;
			12'd152: q <= 1'b1;
			12'd153: q <= 1'b1;
			12'd154: q <= 1'b1;
			12'd155: q <= 1'b1;
			12'd156: q <= 1'b1;
			12'd157: q <= 1'b1;
			12'd158: q <= 1'b1;
			12'd159: q <= 1'b1;
			12'd160: q <= 1'b1;
			12'd161: q <= 1'b1;
			12'd162: q <= 1'b1;
			12'd163: q <= 1'b1;
			12'd164: q <= 1'b1;
			12'd165: q <= 1'b1;
			12'd166: q <= 1'b1;
			12'd167: q <= 1'b1;
			12'd168: q <= 1'b1;
			12'd169: q <= 1'b1;
			12'd170: q <= 1'b1;
			12'd171: q <= 1'b1;
			12'd172: q <= 1'b1;
			12'd173: q <= 1'b1;
			12'd174: q <= 1'b1;
			12'd175: q <= 1'b1;
			12'd176: q <= 1'b1;
			12'd177: q <= 1'b1;
			12'd178: q <= 1'b1;
			12'd179: q <= 1'b1;
			12'd180: q <= 1'b1;
			12'd181: q <= 1'b1;
			12'd182: q <= 1'b1;
			12'd183: q <= 1'b1;
			12'd184: q <= 1'b1;
			12'd185: q <= 1'b1;
			12'd186: q <= 1'b1;
			12'd187: q <= 1'b1;
			12'd188: q <= 1'b1;
			12'd189: q <= 1'b1;
			12'd190: q <= 1'b1;
			12'd191: q <= 1'b1;
			12'd192: q <= 1'b1;
			12'd193: q <= 1'b1;
			12'd194: q <= 1'b1;
			12'd195: q <= 1'b1;
			12'd196: q <= 1'b1;
			12'd197: q <= 1'b1;
			12'd198: q <= 1'b1;
			12'd199: q <= 1'b1;
			12'd200: q <= 1'b1;
			12'd201: q <= 1'b1;
			12'd202: q <= 1'b1;
			12'd203: q <= 1'b1;
			12'd204: q <= 1'b1;
			12'd205: q <= 1'b1;
			12'd206: q <= 1'b1;
			12'd207: q <= 1'b1;
			12'd208: q <= 1'b1;
			12'd209: q <= 1'b1;
			12'd210: q <= 1'b1;
			12'd211: q <= 1'b1;
			12'd212: q <= 1'b1;
			12'd213: q <= 1'b1;
			12'd214: q <= 1'b1;
			12'd215: q <= 1'b1;
			12'd216: q <= 1'b1;
			12'd217: q <= 1'b1;
			12'd218: q <= 1'b1;
			12'd219: q <= 1'b1;
			12'd220: q <= 1'b1;
			12'd221: q <= 1'b1;
			12'd222: q <= 1'b1;
			12'd223: q <= 1'b1;
			12'd224: q <= 1'b1;
			12'd225: q <= 1'b1;
			12'd226: q <= 1'b1;
			12'd227: q <= 1'b1;
			12'd228: q <= 1'b1;
			12'd229: q <= 1'b1;
			12'd230: q <= 1'b1;
			12'd231: q <= 1'b1;
			12'd232: q <= 1'b1;
			12'd233: q <= 1'b1;
			12'd234: q <= 1'b1;
			12'd235: q <= 1'b1;
			12'd236: q <= 1'b1;
			12'd237: q <= 1'b1;
			12'd238: q <= 1'b1;
			12'd239: q <= 1'b1;
			12'd240: q <= 1'b1;
			12'd241: q <= 1'b1;
			12'd242: q <= 1'b1;
			12'd243: q <= 1'b1;
			12'd244: q <= 1'b1;
			12'd245: q <= 1'b1;
			12'd246: q <= 1'b1;
			12'd247: q <= 1'b1;
			12'd248: q <= 1'b1;
			12'd249: q <= 1'b1;
			12'd250: q <= 1'b1;
			12'd251: q <= 1'b1;
			12'd252: q <= 1'b1;
			12'd253: q <= 1'b1;
			12'd254: q <= 1'b1;
			12'd255: q <= 1'b1;
			12'd256: q <= 1'b1;
			12'd257: q <= 1'b1;
			12'd258: q <= 1'b1;
			12'd259: q <= 1'b1;
			12'd260: q <= 1'b1;
			12'd261: q <= 1'b1;
			12'd262: q <= 1'b1;
			12'd263: q <= 1'b1;
			12'd264: q <= 1'b1;
			12'd265: q <= 1'b1;
			12'd266: q <= 1'b1;
			12'd267: q <= 1'b1;
			12'd268: q <= 1'b1;
			12'd269: q <= 1'b1;
			12'd270: q <= 1'b1;
			12'd271: q <= 1'b1;
			12'd272: q <= 1'b1;
			12'd273: q <= 1'b1;
			12'd274: q <= 1'b1;
			12'd275: q <= 1'b1;
			12'd276: q <= 1'b1;
			12'd277: q <= 1'b1;
			12'd278: q <= 1'b1;
			12'd279: q <= 1'b1;
			12'd280: q <= 1'b1;
			12'd281: q <= 1'b1;
			12'd282: q <= 1'b1;
			12'd283: q <= 1'b1;
			12'd284: q <= 1'b1;
			12'd285: q <= 1'b1;
			12'd286: q <= 1'b1;
			12'd287: q <= 1'b1;
			12'd288: q <= 1'b1;
			12'd289: q <= 1'b1;
			12'd290: q <= 1'b1;
			12'd291: q <= 1'b1;
			12'd292: q <= 1'b1;
			12'd293: q <= 1'b1;
			12'd294: q <= 1'b1;
			12'd295: q <= 1'b1;
			12'd296: q <= 1'b1;
			12'd297: q <= 1'b1;
			12'd298: q <= 1'b0;
			12'd299: q <= 1'b0;
			12'd300: q <= 1'b0;
			12'd301: q <= 1'b0;
			12'd302: q <= 1'b1;
			12'd303: q <= 1'b1;
			12'd304: q <= 1'b1;
			12'd305: q <= 1'b1;
			12'd306: q <= 1'b1;
			12'd307: q <= 1'b1;
			12'd308: q <= 1'b1;
			12'd309: q <= 1'b1;
			12'd310: q <= 1'b1;
			12'd311: q <= 1'b1;
			12'd312: q <= 1'b1;
			12'd313: q <= 1'b1;
			12'd314: q <= 1'b1;
			12'd315: q <= 1'b1;
			12'd316: q <= 1'b1;
			12'd317: q <= 1'b1;
			12'd318: q <= 1'b1;
			12'd319: q <= 1'b1;
			12'd320: q <= 1'b1;
			12'd321: q <= 1'b1;
			12'd322: q <= 1'b1;
			12'd323: q <= 1'b1;
			12'd324: q <= 1'b1;
			12'd325: q <= 1'b1;
			12'd326: q <= 1'b1;
			12'd327: q <= 1'b1;
			12'd328: q <= 1'b1;
			12'd329: q <= 1'b1;
			12'd330: q <= 1'b1;
			12'd331: q <= 1'b1;
			12'd332: q <= 1'b1;
			12'd333: q <= 1'b1;
			12'd334: q <= 1'b1;
			12'd335: q <= 1'b1;
			12'd336: q <= 1'b1;
			12'd337: q <= 1'b1;
			12'd338: q <= 1'b1;
			12'd339: q <= 1'b0;
			12'd340: q <= 1'b0;
			12'd341: q <= 1'b0;
			12'd342: q <= 1'b1;
			12'd343: q <= 1'b1;
			12'd344: q <= 1'b1;
			12'd345: q <= 1'b1;
			12'd346: q <= 1'b1;
			12'd347: q <= 1'b1;
			12'd348: q <= 1'b1;
			12'd349: q <= 1'b1;
			12'd350: q <= 1'b1;
			12'd351: q <= 1'b1;
			12'd352: q <= 1'b1;
			12'd353: q <= 1'b1;
			12'd354: q <= 1'b1;
			12'd355: q <= 1'b1;
			12'd356: q <= 1'b1;
			12'd357: q <= 1'b1;
			12'd358: q <= 1'b1;
			12'd359: q <= 1'b1;
			12'd360: q <= 1'b1;
			12'd361: q <= 1'b1;
			12'd362: q <= 1'b1;
			12'd363: q <= 1'b1;
			12'd364: q <= 1'b1;
			12'd365: q <= 1'b1;
			12'd366: q <= 1'b1;
			12'd367: q <= 1'b1;
			12'd368: q <= 1'b1;
			12'd369: q <= 1'b1;
			12'd370: q <= 1'b1;
			12'd371: q <= 1'b1;
			12'd372: q <= 1'b1;
			12'd373: q <= 1'b1;
			12'd374: q <= 1'b1;
			12'd375: q <= 1'b1;
			12'd376: q <= 1'b1;
			12'd377: q <= 1'b1;
			12'd378: q <= 1'b1;
			12'd379: q <= 1'b1;
			12'd380: q <= 1'b1;
			12'd381: q <= 1'b0;
			12'd382: q <= 1'b0;
			12'd383: q <= 1'b0;
			12'd384: q <= 1'b1;
			12'd385: q <= 1'b1;
			12'd386: q <= 1'b1;
			12'd387: q <= 1'b1;
			12'd388: q <= 1'b1;
			12'd389: q <= 1'b1;
			12'd390: q <= 1'b1;
			12'd391: q <= 1'b1;
			12'd392: q <= 1'b1;
			12'd393: q <= 1'b1;
			12'd394: q <= 1'b1;
			12'd395: q <= 1'b1;
			12'd396: q <= 1'b1;
			12'd397: q <= 1'b1;
			12'd398: q <= 1'b1;
			12'd399: q <= 1'b1;
			12'd400: q <= 1'b1;
			12'd401: q <= 1'b1;
			12'd402: q <= 1'b1;
			12'd403: q <= 1'b1;
			12'd404: q <= 1'b1;
			12'd405: q <= 1'b1;
			12'd406: q <= 1'b1;
			12'd407: q <= 1'b1;
			12'd408: q <= 1'b1;
			12'd409: q <= 1'b1;
			12'd410: q <= 1'b1;
			12'd411: q <= 1'b1;
			12'd412: q <= 1'b1;
			12'd413: q <= 1'b1;
			12'd414: q <= 1'b1;
			12'd415: q <= 1'b1;
			12'd416: q <= 1'b1;
			12'd417: q <= 1'b1;
			12'd418: q <= 1'b1;
			12'd419: q <= 1'b1;
			12'd420: q <= 1'b1;
			12'd421: q <= 1'b1;
			12'd422: q <= 1'b1;
			12'd423: q <= 1'b0;
			12'd424: q <= 1'b0;
			12'd425: q <= 1'b1;
			12'd426: q <= 1'b1;
			12'd427: q <= 1'b1;
			12'd428: q <= 1'b1;
			12'd429: q <= 1'b1;
			12'd430: q <= 1'b1;
			12'd431: q <= 1'b1;
			12'd432: q <= 1'b1;
			12'd433: q <= 1'b1;
			12'd434: q <= 1'b1;
			12'd435: q <= 1'b1;
			12'd436: q <= 1'b1;
			12'd437: q <= 1'b1;
			12'd438: q <= 1'b1;
			12'd439: q <= 1'b1;
			12'd440: q <= 1'b1;
			12'd441: q <= 1'b1;
			12'd442: q <= 1'b1;
			12'd443: q <= 1'b1;
			12'd444: q <= 1'b1;
			12'd445: q <= 1'b1;
			12'd446: q <= 1'b1;
			12'd447: q <= 1'b1;
			12'd448: q <= 1'b1;
			12'd449: q <= 1'b1;
			12'd450: q <= 1'b1;
			12'd451: q <= 1'b1;
			12'd452: q <= 1'b1;
			12'd453: q <= 1'b1;
			12'd454: q <= 1'b1;
			12'd455: q <= 1'b1;
			12'd456: q <= 1'b1;
			12'd457: q <= 1'b1;
			12'd458: q <= 1'b1;
			12'd459: q <= 1'b1;
			12'd460: q <= 1'b1;
			12'd461: q <= 1'b1;
			12'd462: q <= 1'b1;
			12'd463: q <= 1'b1;
			12'd464: q <= 1'b1;
			12'd465: q <= 1'b0;
			12'd466: q <= 1'b0;
			12'd467: q <= 1'b1;
			12'd468: q <= 1'b1;
			12'd469: q <= 1'b1;
			12'd470: q <= 1'b1;
			12'd471: q <= 1'b1;
			12'd472: q <= 1'b1;
			12'd473: q <= 1'b1;
			12'd474: q <= 1'b1;
			12'd475: q <= 1'b1;
			12'd476: q <= 1'b1;
			12'd477: q <= 1'b1;
			12'd478: q <= 1'b1;
			12'd479: q <= 1'b1;
			12'd480: q <= 1'b1;
			12'd481: q <= 1'b1;
			12'd482: q <= 1'b1;
			12'd483: q <= 1'b1;
			12'd484: q <= 1'b1;
			12'd485: q <= 1'b1;
			12'd486: q <= 1'b1;
			12'd487: q <= 1'b1;
			12'd488: q <= 1'b1;
			12'd489: q <= 1'b1;
			12'd490: q <= 1'b1;
			12'd491: q <= 1'b1;
			12'd492: q <= 1'b1;
			12'd493: q <= 1'b1;
			12'd494: q <= 1'b1;
			12'd495: q <= 1'b1;
			12'd496: q <= 1'b1;
			12'd497: q <= 1'b1;
			12'd498: q <= 1'b1;
			12'd499: q <= 1'b1;
			12'd500: q <= 1'b1;
			12'd501: q <= 1'b1;
			12'd502: q <= 1'b1;
			12'd503: q <= 1'b1;
			12'd504: q <= 1'b1;
			12'd505: q <= 1'b1;
			12'd506: q <= 1'b0;
			12'd507: q <= 1'b0;
			12'd508: q <= 1'b0;
			12'd509: q <= 1'b0;
			12'd510: q <= 1'b1;
			12'd511: q <= 1'b1;
			12'd512: q <= 1'b1;
			12'd513: q <= 1'b1;
			12'd514: q <= 1'b1;
			12'd515: q <= 1'b1;
			12'd516: q <= 1'b1;
			12'd517: q <= 1'b1;
			12'd518: q <= 1'b1;
			12'd519: q <= 1'b1;
			12'd520: q <= 1'b1;
			12'd521: q <= 1'b1;
			12'd522: q <= 1'b1;
			12'd523: q <= 1'b1;
			12'd524: q <= 1'b1;
			12'd525: q <= 1'b1;
			12'd526: q <= 1'b1;
			12'd527: q <= 1'b1;
			12'd528: q <= 1'b1;
			12'd529: q <= 1'b1;
			12'd530: q <= 1'b1;
			12'd531: q <= 1'b1;
			12'd532: q <= 1'b1;
			12'd533: q <= 1'b1;
			12'd534: q <= 1'b1;
			12'd535: q <= 1'b1;
			12'd536: q <= 1'b1;
			12'd537: q <= 1'b1;
			12'd538: q <= 1'b1;
			12'd539: q <= 1'b1;
			12'd540: q <= 1'b1;
			12'd541: q <= 1'b1;
			12'd542: q <= 1'b1;
			12'd543: q <= 1'b1;
			12'd544: q <= 1'b1;
			12'd545: q <= 1'b1;
			12'd546: q <= 1'b1;
			12'd547: q <= 1'b1;
			12'd548: q <= 1'b1;
			12'd549: q <= 1'b1;
			12'd550: q <= 1'b1;
			12'd551: q <= 1'b1;
			12'd552: q <= 1'b1;
			12'd553: q <= 1'b1;
			12'd554: q <= 1'b1;
			12'd555: q <= 1'b1;
			12'd556: q <= 1'b1;
			12'd557: q <= 1'b1;
			12'd558: q <= 1'b1;
			12'd559: q <= 1'b1;
			12'd560: q <= 1'b1;
			12'd561: q <= 1'b1;
			12'd562: q <= 1'b1;
			12'd563: q <= 1'b1;
			12'd564: q <= 1'b1;
			12'd565: q <= 1'b1;
			12'd566: q <= 1'b1;
			12'd567: q <= 1'b1;
			12'd568: q <= 1'b1;
			12'd569: q <= 1'b1;
			12'd570: q <= 1'b1;
			12'd571: q <= 1'b1;
			12'd572: q <= 1'b1;
			12'd573: q <= 1'b1;
			12'd574: q <= 1'b1;
			12'd575: q <= 1'b1;
			12'd576: q <= 1'b1;
			12'd577: q <= 1'b1;
			12'd578: q <= 1'b1;
			12'd579: q <= 1'b1;
			12'd580: q <= 1'b1;
			12'd581: q <= 1'b1;
			12'd582: q <= 1'b1;
			12'd583: q <= 1'b1;
			12'd584: q <= 1'b1;
			12'd585: q <= 1'b1;
			12'd586: q <= 1'b1;
			12'd587: q <= 1'b1;
			12'd588: q <= 1'b1;
			12'd589: q <= 1'b1;
			12'd590: q <= 1'b1;
			12'd591: q <= 1'b1;
			12'd592: q <= 1'b1;
			12'd593: q <= 1'b1;
			12'd594: q <= 1'b1;
			12'd595: q <= 1'b1;
			12'd596: q <= 1'b1;
			12'd597: q <= 1'b1;
			12'd598: q <= 1'b1;
			12'd599: q <= 1'b1;
			12'd600: q <= 1'b1;
			12'd601: q <= 1'b1;
			12'd602: q <= 1'b1;
			12'd603: q <= 1'b1;
			12'd604: q <= 1'b1;
			12'd605: q <= 1'b1;
			12'd606: q <= 1'b1;
			12'd607: q <= 1'b1;
			12'd608: q <= 1'b1;
			12'd609: q <= 1'b1;
			12'd610: q <= 1'b1;
			12'd611: q <= 1'b1;
			12'd612: q <= 1'b0;
			12'd613: q <= 1'b0;
			12'd614: q <= 1'b0;
			12'd615: q <= 1'b0;
			12'd616: q <= 1'b1;
			12'd617: q <= 1'b1;
			12'd618: q <= 1'b1;
			12'd619: q <= 1'b1;
			12'd620: q <= 1'b1;
			12'd621: q <= 1'b1;
			12'd622: q <= 1'b1;
			12'd623: q <= 1'b1;
			12'd624: q <= 1'b1;
			12'd625: q <= 1'b1;
			12'd626: q <= 1'b0;
			12'd627: q <= 1'b0;
			12'd628: q <= 1'b0;
			12'd629: q <= 1'b0;
			12'd630: q <= 1'b0;
			12'd631: q <= 1'b1;
			12'd632: q <= 1'b1;
			12'd633: q <= 1'b1;
			12'd634: q <= 1'b1;
			12'd635: q <= 1'b1;
			12'd636: q <= 1'b1;
			12'd637: q <= 1'b1;
			12'd638: q <= 1'b1;
			12'd639: q <= 1'b1;
			12'd640: q <= 1'b1;
			12'd641: q <= 1'b1;
			12'd642: q <= 1'b1;
			12'd643: q <= 1'b1;
			12'd644: q <= 1'b1;
			12'd645: q <= 1'b1;
			12'd646: q <= 1'b1;
			12'd647: q <= 1'b1;
			12'd648: q <= 1'b1;
			12'd649: q <= 1'b1;
			12'd650: q <= 1'b0;
			12'd651: q <= 1'b0;
			12'd652: q <= 1'b0;
			12'd653: q <= 1'b0;
			12'd654: q <= 1'b0;
			12'd655: q <= 1'b0;
			12'd656: q <= 1'b0;
			12'd657: q <= 1'b0;
			12'd658: q <= 1'b1;
			12'd659: q <= 1'b1;
			12'd660: q <= 1'b1;
			12'd661: q <= 1'b1;
			12'd662: q <= 1'b1;
			12'd663: q <= 1'b1;
			12'd664: q <= 1'b0;
			12'd665: q <= 1'b0;
			12'd666: q <= 1'b0;
			12'd667: q <= 1'b0;
			12'd668: q <= 1'b0;
			12'd669: q <= 1'b0;
			12'd670: q <= 1'b0;
			12'd671: q <= 1'b0;
			12'd672: q <= 1'b0;
			12'd673: q <= 1'b0;
			12'd674: q <= 1'b1;
			12'd675: q <= 1'b1;
			12'd676: q <= 1'b1;
			12'd677: q <= 1'b1;
			12'd678: q <= 1'b1;
			12'd679: q <= 1'b1;
			12'd680: q <= 1'b1;
			12'd681: q <= 1'b1;
			12'd682: q <= 1'b1;
			12'd683: q <= 1'b1;
			12'd684: q <= 1'b1;
			12'd685: q <= 1'b1;
			12'd686: q <= 1'b1;
			12'd687: q <= 1'b1;
			12'd688: q <= 1'b1;
			12'd689: q <= 1'b0;
			12'd690: q <= 1'b0;
			12'd691: q <= 1'b0;
			12'd692: q <= 1'b0;
			12'd693: q <= 1'b0;
			12'd694: q <= 1'b0;
			12'd695: q <= 1'b0;
			12'd696: q <= 1'b0;
			12'd697: q <= 1'b0;
			12'd698: q <= 1'b0;
			12'd699: q <= 1'b0;
			12'd700: q <= 1'b1;
			12'd701: q <= 1'b1;
			12'd702: q <= 1'b1;
			12'd703: q <= 1'b1;
			12'd704: q <= 1'b1;
			12'd705: q <= 1'b1;
			12'd706: q <= 1'b0;
			12'd707: q <= 1'b0;
			12'd708: q <= 1'b0;
			12'd709: q <= 1'b0;
			12'd710: q <= 1'b0;
			12'd711: q <= 1'b0;
			12'd712: q <= 1'b0;
			12'd713: q <= 1'b0;
			12'd714: q <= 1'b0;
			12'd715: q <= 1'b1;
			12'd716: q <= 1'b1;
			12'd717: q <= 1'b1;
			12'd718: q <= 1'b1;
			12'd719: q <= 1'b1;
			12'd720: q <= 1'b1;
			12'd721: q <= 1'b1;
			12'd722: q <= 1'b1;
			12'd723: q <= 1'b1;
			12'd724: q <= 1'b1;
			12'd725: q <= 1'b1;
			12'd726: q <= 1'b1;
			12'd727: q <= 1'b1;
			12'd728: q <= 1'b1;
			12'd729: q <= 1'b0;
			12'd730: q <= 1'b0;
			12'd731: q <= 1'b0;
			12'd732: q <= 1'b0;
			12'd733: q <= 1'b0;
			12'd734: q <= 1'b0;
			12'd735: q <= 1'b0;
			12'd736: q <= 1'b0;
			12'd737: q <= 1'b0;
			12'd738: q <= 1'b0;
			12'd739: q <= 1'b0;
			12'd740: q <= 1'b0;
			12'd741: q <= 1'b1;
			12'd742: q <= 1'b1;
			12'd743: q <= 1'b1;
			12'd744: q <= 1'b1;
			12'd745: q <= 1'b1;
			12'd746: q <= 1'b0;
			12'd747: q <= 1'b0;
			12'd748: q <= 1'b0;
			12'd749: q <= 1'b0;
			12'd750: q <= 1'b0;
			12'd751: q <= 1'b0;
			12'd752: q <= 1'b0;
			12'd753: q <= 1'b0;
			12'd754: q <= 1'b0;
			12'd755: q <= 1'b1;
			12'd756: q <= 1'b1;
			12'd757: q <= 1'b1;
			12'd758: q <= 1'b1;
			12'd759: q <= 1'b1;
			12'd760: q <= 1'b1;
			12'd761: q <= 1'b1;
			12'd762: q <= 1'b1;
			12'd763: q <= 1'b1;
			12'd764: q <= 1'b1;
			12'd765: q <= 1'b1;
			12'd766: q <= 1'b1;
			12'd767: q <= 1'b1;
			12'd768: q <= 1'b0;
			12'd769: q <= 1'b0;
			12'd770: q <= 1'b0;
			12'd771: q <= 1'b0;
			12'd772: q <= 1'b0;
			12'd773: q <= 1'b0;
			12'd774: q <= 1'b0;
			12'd775: q <= 1'b0;
			12'd776: q <= 1'b0;
			12'd777: q <= 1'b0;
			12'd778: q <= 1'b0;
			12'd779: q <= 1'b0;
			12'd780: q <= 1'b0;
			12'd781: q <= 1'b1;
			12'd782: q <= 1'b1;
			12'd783: q <= 1'b1;
			12'd784: q <= 1'b1;
			12'd785: q <= 1'b1;
			12'd786: q <= 1'b0;
			12'd787: q <= 1'b0;
			12'd788: q <= 1'b0;
			12'd789: q <= 1'b0;
			12'd790: q <= 1'b0;
			12'd791: q <= 1'b0;
			12'd792: q <= 1'b0;
			12'd793: q <= 1'b0;
			12'd794: q <= 1'b0;
			12'd795: q <= 1'b0;
			12'd796: q <= 1'b1;
			12'd797: q <= 1'b1;
			12'd798: q <= 1'b1;
			12'd799: q <= 1'b1;
			12'd800: q <= 1'b1;
			12'd801: q <= 1'b1;
			12'd802: q <= 1'b1;
			12'd803: q <= 1'b1;
			12'd804: q <= 1'b1;
			12'd805: q <= 1'b1;
			12'd806: q <= 1'b1;
			12'd807: q <= 1'b1;
			12'd808: q <= 1'b1;
			12'd809: q <= 1'b0;
			12'd810: q <= 1'b0;
			12'd811: q <= 1'b0;
			12'd812: q <= 1'b0;
			12'd813: q <= 1'b0;
			12'd814: q <= 1'b0;
			12'd815: q <= 1'b0;
			12'd816: q <= 1'b0;
			12'd817: q <= 1'b0;
			12'd818: q <= 1'b0;
			12'd819: q <= 1'b0;
			12'd820: q <= 1'b0;
			12'd821: q <= 1'b0;
			12'd822: q <= 1'b1;
			12'd823: q <= 1'b1;
			12'd824: q <= 1'b1;
			12'd825: q <= 1'b1;
			12'd826: q <= 1'b1;
			12'd827: q <= 1'b0;
			12'd828: q <= 1'b0;
			12'd829: q <= 1'b0;
			12'd830: q <= 1'b0;
			12'd831: q <= 1'b0;
			12'd832: q <= 1'b0;
			12'd833: q <= 1'b0;
			12'd834: q <= 1'b0;
			12'd835: q <= 1'b0;
			12'd836: q <= 1'b1;
			12'd837: q <= 1'b1;
			12'd838: q <= 1'b1;
			12'd839: q <= 1'b1;
			12'd840: q <= 1'b1;
			12'd841: q <= 1'b1;
			12'd842: q <= 1'b1;
			12'd843: q <= 1'b1;
			12'd844: q <= 1'b1;
			12'd845: q <= 1'b1;
			12'd846: q <= 1'b1;
			12'd847: q <= 1'b1;
			12'd848: q <= 1'b1;
			12'd849: q <= 1'b0;
			12'd850: q <= 1'b0;
			12'd851: q <= 1'b0;
			12'd852: q <= 1'b0;
			12'd853: q <= 1'b0;
			12'd854: q <= 1'b0;
			12'd855: q <= 1'b0;
			12'd856: q <= 1'b0;
			12'd857: q <= 1'b0;
			12'd858: q <= 1'b0;
			12'd859: q <= 1'b0;
			12'd860: q <= 1'b0;
			12'd861: q <= 1'b0;
			12'd862: q <= 1'b1;
			12'd863: q <= 1'b1;
			12'd864: q <= 1'b1;
			12'd865: q <= 1'b1;
			12'd866: q <= 1'b1;
			12'd867: q <= 1'b0;
			12'd868: q <= 1'b0;
			12'd869: q <= 1'b0;
			12'd870: q <= 1'b0;
			12'd871: q <= 1'b0;
			12'd872: q <= 1'b0;
			12'd873: q <= 1'b0;
			12'd874: q <= 1'b0;
			12'd875: q <= 1'b1;
			12'd876: q <= 1'b1;
			12'd877: q <= 1'b1;
			12'd878: q <= 1'b1;
			12'd879: q <= 1'b1;
			12'd880: q <= 1'b1;
			12'd881: q <= 1'b1;
			12'd882: q <= 1'b1;
			12'd883: q <= 1'b1;
			12'd884: q <= 1'b1;
			12'd885: q <= 1'b1;
			12'd886: q <= 1'b1;
			12'd887: q <= 1'b1;
			12'd888: q <= 1'b1;
			12'd889: q <= 1'b0;
			12'd890: q <= 1'b0;
			12'd891: q <= 1'b0;
			12'd892: q <= 1'b0;
			12'd893: q <= 1'b0;
			12'd894: q <= 1'b0;
			12'd895: q <= 1'b0;
			12'd896: q <= 1'b0;
			12'd897: q <= 1'b0;
			12'd898: q <= 1'b0;
			12'd899: q <= 1'b0;
			12'd900: q <= 1'b0;
			12'd901: q <= 1'b0;
			12'd902: q <= 1'b1;
			12'd903: q <= 1'b1;
			12'd904: q <= 1'b1;
			12'd905: q <= 1'b1;
			12'd906: q <= 1'b1;
			12'd907: q <= 1'b0;
			12'd908: q <= 1'b0;
			12'd909: q <= 1'b0;
			12'd910: q <= 1'b0;
			12'd911: q <= 1'b0;
			12'd912: q <= 1'b0;
			12'd913: q <= 1'b0;
			12'd914: q <= 1'b0;
			12'd915: q <= 1'b1;
			12'd916: q <= 1'b1;
			12'd917: q <= 1'b1;
			12'd918: q <= 1'b1;
			12'd919: q <= 1'b1;
			12'd920: q <= 1'b1;
			12'd921: q <= 1'b1;
			12'd922: q <= 1'b1;
			12'd923: q <= 1'b1;
			12'd924: q <= 1'b1;
			12'd925: q <= 1'b1;
			12'd926: q <= 1'b1;
			12'd927: q <= 1'b1;
			12'd928: q <= 1'b0;
			12'd929: q <= 1'b0;
			12'd930: q <= 1'b0;
			12'd931: q <= 1'b0;
			12'd932: q <= 1'b0;
			12'd933: q <= 1'b0;
			12'd934: q <= 1'b0;
			12'd935: q <= 1'b0;
			12'd936: q <= 1'b0;
			12'd937: q <= 1'b0;
			12'd938: q <= 1'b0;
			12'd939: q <= 1'b0;
			12'd940: q <= 1'b0;
			12'd941: q <= 1'b0;
			12'd942: q <= 1'b1;
			12'd943: q <= 1'b1;
			12'd944: q <= 1'b1;
			12'd945: q <= 1'b1;
			12'd946: q <= 1'b1;
			12'd947: q <= 1'b0;
			12'd948: q <= 1'b0;
			12'd949: q <= 1'b0;
			12'd950: q <= 1'b0;
			12'd951: q <= 1'b0;
			12'd952: q <= 1'b0;
			12'd953: q <= 1'b0;
			12'd954: q <= 1'b0;
			12'd955: q <= 1'b1;
			12'd956: q <= 1'b1;
			12'd957: q <= 1'b1;
			12'd958: q <= 1'b1;
			12'd959: q <= 1'b1;
			12'd960: q <= 1'b1;
			12'd961: q <= 1'b1;
			12'd962: q <= 1'b1;
			12'd963: q <= 1'b1;
			12'd964: q <= 1'b1;
			12'd965: q <= 1'b1;
			12'd966: q <= 1'b1;
			12'd967: q <= 1'b1;
			12'd968: q <= 1'b0;
			12'd969: q <= 1'b0;
			12'd970: q <= 1'b0;
			12'd971: q <= 1'b0;
			12'd972: q <= 1'b0;
			12'd973: q <= 1'b0;
			12'd974: q <= 1'b0;
			12'd975: q <= 1'b0;
			12'd976: q <= 1'b0;
			12'd977: q <= 1'b0;
			12'd978: q <= 1'b0;
			12'd979: q <= 1'b0;
			12'd980: q <= 1'b0;
			12'd981: q <= 1'b0;
			12'd982: q <= 1'b0;
			12'd983: q <= 1'b1;
			12'd984: q <= 1'b1;
			12'd985: q <= 1'b1;
			12'd986: q <= 1'b0;
			12'd987: q <= 1'b0;
			12'd988: q <= 1'b0;
			12'd989: q <= 1'b0;
			12'd990: q <= 1'b0;
			12'd991: q <= 1'b0;
			12'd992: q <= 1'b0;
			12'd993: q <= 1'b0;
			12'd994: q <= 1'b1;
			12'd995: q <= 1'b1;
			12'd996: q <= 1'b1;
			12'd997: q <= 1'b1;
			12'd998: q <= 1'b1;
			12'd999: q <= 1'b1;
			12'd1000: q <= 1'b1;
			12'd1001: q <= 1'b1;
			12'd1002: q <= 1'b1;
			12'd1003: q <= 1'b1;
			12'd1004: q <= 1'b1;
			12'd1005: q <= 1'b1;
			12'd1006: q <= 1'b1;
			12'd1007: q <= 1'b1;
			12'd1008: q <= 1'b0;
			12'd1009: q <= 1'b0;
			12'd1010: q <= 1'b0;
			12'd1011: q <= 1'b0;
			12'd1012: q <= 1'b0;
			12'd1013: q <= 1'b0;
			12'd1014: q <= 1'b0;
			12'd1015: q <= 1'b0;
			12'd1016: q <= 1'b0;
			12'd1017: q <= 1'b0;
			12'd1018: q <= 1'b0;
			12'd1019: q <= 1'b0;
			12'd1020: q <= 1'b0;
			12'd1021: q <= 1'b0;
			12'd1022: q <= 1'b0;
			12'd1023: q <= 1'b0;
			12'd1024: q <= 1'b0;
			12'd1025: q <= 1'b0;
			12'd1026: q <= 1'b0;
			12'd1027: q <= 1'b0;
			12'd1028: q <= 1'b0;
			12'd1029: q <= 1'b0;
			12'd1030: q <= 1'b0;
			12'd1031: q <= 1'b0;
			12'd1032: q <= 1'b0;
			12'd1033: q <= 1'b0;
			12'd1034: q <= 1'b1;
			12'd1035: q <= 1'b1;
			12'd1036: q <= 1'b1;
			12'd1037: q <= 1'b1;
			12'd1038: q <= 1'b1;
			12'd1039: q <= 1'b1;
			12'd1040: q <= 1'b1;
			12'd1041: q <= 1'b1;
			12'd1042: q <= 1'b1;
			12'd1043: q <= 1'b1;
			12'd1044: q <= 1'b1;
			12'd1045: q <= 1'b1;
			12'd1046: q <= 1'b1;
			12'd1047: q <= 1'b1;
			12'd1048: q <= 1'b0;
			12'd1049: q <= 1'b0;
			12'd1050: q <= 1'b0;
			12'd1051: q <= 1'b0;
			12'd1052: q <= 1'b0;
			12'd1053: q <= 1'b0;
			12'd1054: q <= 1'b0;
			12'd1055: q <= 1'b0;
			12'd1056: q <= 1'b0;
			12'd1057: q <= 1'b0;
			12'd1058: q <= 1'b0;
			12'd1059: q <= 1'b0;
			12'd1060: q <= 1'b0;
			12'd1061: q <= 1'b0;
			12'd1062: q <= 1'b0;
			12'd1063: q <= 1'b0;
			12'd1064: q <= 1'b0;
			12'd1065: q <= 1'b0;
			12'd1066: q <= 1'b0;
			12'd1067: q <= 1'b0;
			12'd1068: q <= 1'b0;
			12'd1069: q <= 1'b0;
			12'd1070: q <= 1'b0;
			12'd1071: q <= 1'b0;
			12'd1072: q <= 1'b0;
			12'd1073: q <= 1'b1;
			12'd1074: q <= 1'b1;
			12'd1075: q <= 1'b1;
			12'd1076: q <= 1'b1;
			12'd1077: q <= 1'b1;
			12'd1078: q <= 1'b1;
			12'd1079: q <= 1'b1;
			12'd1080: q <= 1'b1;
			12'd1081: q <= 1'b1;
			12'd1082: q <= 1'b1;
			12'd1083: q <= 1'b1;
			12'd1084: q <= 1'b1;
			12'd1085: q <= 1'b1;
			12'd1086: q <= 1'b1;
			12'd1087: q <= 1'b1;
			12'd1088: q <= 1'b0;
			12'd1089: q <= 1'b0;
			12'd1090: q <= 1'b0;
			12'd1091: q <= 1'b0;
			12'd1092: q <= 1'b0;
			12'd1093: q <= 1'b0;
			12'd1094: q <= 1'b0;
			12'd1095: q <= 1'b0;
			12'd1096: q <= 1'b0;
			12'd1097: q <= 1'b0;
			12'd1098: q <= 1'b0;
			12'd1099: q <= 1'b0;
			12'd1100: q <= 1'b0;
			12'd1101: q <= 1'b0;
			12'd1102: q <= 1'b0;
			12'd1103: q <= 1'b0;
			12'd1104: q <= 1'b0;
			12'd1105: q <= 1'b0;
			12'd1106: q <= 1'b0;
			12'd1107: q <= 1'b0;
			12'd1108: q <= 1'b0;
			12'd1109: q <= 1'b0;
			12'd1110: q <= 1'b0;
			12'd1111: q <= 1'b0;
			12'd1112: q <= 1'b0;
			12'd1113: q <= 1'b1;
			12'd1114: q <= 1'b1;
			12'd1115: q <= 1'b1;
			12'd1116: q <= 1'b1;
			12'd1117: q <= 1'b1;
			12'd1118: q <= 1'b1;
			12'd1119: q <= 1'b1;
			12'd1120: q <= 1'b0;
			12'd1121: q <= 1'b0;
			12'd1122: q <= 1'b0;
			12'd1123: q <= 1'b0;
			12'd1124: q <= 1'b0;
			12'd1125: q <= 1'b0;
			12'd1126: q <= 1'b0;
			12'd1127: q <= 1'b0;
			12'd1128: q <= 1'b0;
			12'd1129: q <= 1'b0;
			12'd1130: q <= 1'b0;
			12'd1131: q <= 1'b0;
			12'd1132: q <= 1'b0;
			12'd1133: q <= 1'b0;
			12'd1134: q <= 1'b0;
			12'd1135: q <= 1'b0;
			12'd1136: q <= 1'b0;
			12'd1137: q <= 1'b0;
			12'd1138: q <= 1'b0;
			12'd1139: q <= 1'b0;
			12'd1140: q <= 1'b0;
			12'd1141: q <= 1'b0;
			12'd1142: q <= 1'b0;
			12'd1143: q <= 1'b0;
			12'd1144: q <= 1'b0;
			12'd1145: q <= 1'b0;
			12'd1146: q <= 1'b0;
			12'd1147: q <= 1'b0;
			12'd1148: q <= 1'b0;
			12'd1149: q <= 1'b0;
			12'd1150: q <= 1'b0;
			12'd1151: q <= 1'b0;
			12'd1152: q <= 1'b1;
			12'd1153: q <= 1'b1;
			12'd1154: q <= 1'b1;
			12'd1155: q <= 1'b1;
			12'd1156: q <= 1'b1;
			12'd1157: q <= 1'b1;
			12'd1158: q <= 1'b1;
			12'd1159: q <= 1'b1;
			12'd1160: q <= 1'b0;
			12'd1161: q <= 1'b0;
			12'd1162: q <= 1'b0;
			12'd1163: q <= 1'b0;
			12'd1164: q <= 1'b0;
			12'd1165: q <= 1'b0;
			12'd1166: q <= 1'b0;
			12'd1167: q <= 1'b0;
			12'd1168: q <= 1'b0;
			12'd1169: q <= 1'b0;
			12'd1170: q <= 1'b0;
			12'd1171: q <= 1'b0;
			12'd1172: q <= 1'b0;
			12'd1173: q <= 1'b0;
			12'd1174: q <= 1'b0;
			12'd1175: q <= 1'b0;
			12'd1176: q <= 1'b0;
			12'd1177: q <= 1'b0;
			12'd1178: q <= 1'b0;
			12'd1179: q <= 1'b0;
			12'd1180: q <= 1'b0;
			12'd1181: q <= 1'b0;
			12'd1182: q <= 1'b0;
			12'd1183: q <= 1'b0;
			12'd1184: q <= 1'b0;
			12'd1185: q <= 1'b0;
			12'd1186: q <= 1'b0;
			12'd1187: q <= 1'b0;
			12'd1188: q <= 1'b0;
			12'd1189: q <= 1'b0;
			12'd1190: q <= 1'b0;
			12'd1191: q <= 1'b0;
			12'd1192: q <= 1'b0;
			12'd1193: q <= 1'b0;
			12'd1194: q <= 1'b0;
			12'd1195: q <= 1'b0;
			12'd1196: q <= 1'b0;
			12'd1197: q <= 1'b0;
			12'd1198: q <= 1'b0;
			12'd1199: q <= 1'b0;
			12'd1200: q <= 1'b0;
			12'd1201: q <= 1'b0;
			12'd1202: q <= 1'b0;
			12'd1203: q <= 1'b0;
			12'd1204: q <= 1'b0;
			12'd1205: q <= 1'b0;
			12'd1206: q <= 1'b0;
			12'd1207: q <= 1'b0;
			12'd1208: q <= 1'b0;
			12'd1209: q <= 1'b0;
			12'd1210: q <= 1'b0;
			12'd1211: q <= 1'b0;
			12'd1212: q <= 1'b0;
			12'd1213: q <= 1'b0;
			12'd1214: q <= 1'b0;
			12'd1215: q <= 1'b0;
			12'd1216: q <= 1'b0;
			12'd1217: q <= 1'b0;
			12'd1218: q <= 1'b0;
			12'd1219: q <= 1'b0;
			12'd1220: q <= 1'b0;
			12'd1221: q <= 1'b0;
			12'd1222: q <= 1'b0;
			12'd1223: q <= 1'b0;
			12'd1224: q <= 1'b0;
			12'd1225: q <= 1'b0;
			12'd1226: q <= 1'b0;
			12'd1227: q <= 1'b0;
			12'd1228: q <= 1'b0;
			12'd1229: q <= 1'b0;
			12'd1230: q <= 1'b0;
			12'd1231: q <= 1'b0;
			12'd1232: q <= 1'b0;
			12'd1233: q <= 1'b0;
			12'd1234: q <= 1'b0;
			12'd1235: q <= 1'b0;
			12'd1236: q <= 1'b0;
			12'd1237: q <= 1'b0;
			12'd1238: q <= 1'b0;
			12'd1239: q <= 1'b0;
			12'd1240: q <= 1'b0;
			12'd1241: q <= 1'b0;
			12'd1242: q <= 1'b0;
			12'd1243: q <= 1'b0;
			12'd1244: q <= 1'b0;
			12'd1245: q <= 1'b0;
			12'd1246: q <= 1'b0;
			12'd1247: q <= 1'b0;
			12'd1248: q <= 1'b0;
			12'd1249: q <= 1'b0;
			12'd1250: q <= 1'b0;
			12'd1251: q <= 1'b0;
			12'd1252: q <= 1'b0;
			12'd1253: q <= 1'b0;
			12'd1254: q <= 1'b0;
			12'd1255: q <= 1'b0;
			12'd1256: q <= 1'b0;
			12'd1257: q <= 1'b0;
			12'd1258: q <= 1'b0;
			12'd1259: q <= 1'b0;
			12'd1260: q <= 1'b0;
			12'd1261: q <= 1'b0;
			12'd1262: q <= 1'b0;
			12'd1263: q <= 1'b0;
			12'd1264: q <= 1'b0;
			12'd1265: q <= 1'b0;
			12'd1266: q <= 1'b0;
			12'd1267: q <= 1'b0;
			12'd1268: q <= 1'b0;
			12'd1269: q <= 1'b0;
			12'd1270: q <= 1'b0;
			12'd1271: q <= 1'b0;
			12'd1272: q <= 1'b0;
			12'd1273: q <= 1'b0;
			12'd1274: q <= 1'b0;
			12'd1275: q <= 1'b0;
			12'd1276: q <= 1'b0;
			12'd1277: q <= 1'b0;
			12'd1278: q <= 1'b0;
			12'd1279: q <= 1'b0;
			12'd1280: q <= 1'b1;
			12'd1281: q <= 1'b1;
			12'd1282: q <= 1'b1;
			12'd1283: q <= 1'b1;
			12'd1284: q <= 1'b0;
			12'd1285: q <= 1'b0;
			12'd1286: q <= 1'b0;
			12'd1287: q <= 1'b0;
			12'd1288: q <= 1'b0;
			12'd1289: q <= 1'b0;
			12'd1290: q <= 1'b0;
			12'd1291: q <= 1'b0;
			12'd1292: q <= 1'b0;
			12'd1293: q <= 1'b0;
			12'd1294: q <= 1'b0;
			12'd1295: q <= 1'b0;
			12'd1296: q <= 1'b0;
			12'd1297: q <= 1'b0;
			12'd1298: q <= 1'b0;
			12'd1299: q <= 1'b0;
			12'd1300: q <= 1'b0;
			12'd1301: q <= 1'b0;
			12'd1302: q <= 1'b0;
			12'd1303: q <= 1'b0;
			12'd1304: q <= 1'b0;
			12'd1305: q <= 1'b0;
			12'd1306: q <= 1'b0;
			12'd1307: q <= 1'b0;
			12'd1308: q <= 1'b0;
			12'd1309: q <= 1'b0;
			12'd1310: q <= 1'b0;
			12'd1311: q <= 1'b0;
			12'd1312: q <= 1'b0;
			12'd1313: q <= 1'b0;
			12'd1314: q <= 1'b0;
			12'd1315: q <= 1'b0;
			12'd1316: q <= 1'b0;
			12'd1317: q <= 1'b0;
			12'd1318: q <= 1'b0;
			12'd1319: q <= 1'b0;
			12'd1320: q <= 1'b1;
			12'd1321: q <= 1'b1;
			12'd1322: q <= 1'b1;
			12'd1323: q <= 1'b1;
			12'd1324: q <= 1'b1;
			12'd1325: q <= 1'b1;
			12'd1326: q <= 1'b0;
			12'd1327: q <= 1'b0;
			12'd1328: q <= 1'b0;
			12'd1329: q <= 1'b0;
			12'd1330: q <= 1'b0;
			12'd1331: q <= 1'b0;
			12'd1332: q <= 1'b0;
			12'd1333: q <= 1'b0;
			12'd1334: q <= 1'b0;
			12'd1335: q <= 1'b0;
			12'd1336: q <= 1'b0;
			12'd1337: q <= 1'b0;
			12'd1338: q <= 1'b0;
			12'd1339: q <= 1'b0;
			12'd1340: q <= 1'b0;
			12'd1341: q <= 1'b0;
			12'd1342: q <= 1'b0;
			12'd1343: q <= 1'b0;
			12'd1344: q <= 1'b0;
			12'd1345: q <= 1'b0;
			12'd1346: q <= 1'b0;
			12'd1347: q <= 1'b0;
			12'd1348: q <= 1'b0;
			12'd1349: q <= 1'b0;
			12'd1350: q <= 1'b0;
			12'd1351: q <= 1'b0;
			12'd1352: q <= 1'b0;
			12'd1353: q <= 1'b1;
			12'd1354: q <= 1'b1;
			12'd1355: q <= 1'b1;
			12'd1356: q <= 1'b1;
			12'd1357: q <= 1'b0;
			12'd1358: q <= 1'b1;
			12'd1359: q <= 1'b0;
			12'd1360: q <= 1'b1;
			12'd1361: q <= 1'b1;
			12'd1362: q <= 1'b1;
			12'd1363: q <= 1'b1;
			12'd1364: q <= 1'b1;
			12'd1365: q <= 1'b1;
			12'd1366: q <= 1'b1;
			12'd1367: q <= 1'b0;
			12'd1368: q <= 1'b0;
			12'd1369: q <= 1'b0;
			12'd1370: q <= 1'b0;
			12'd1371: q <= 1'b0;
			12'd1372: q <= 1'b0;
			12'd1373: q <= 1'b0;
			12'd1374: q <= 1'b0;
			12'd1375: q <= 1'b0;
			12'd1376: q <= 1'b0;
			12'd1377: q <= 1'b0;
			12'd1378: q <= 1'b0;
			12'd1379: q <= 1'b0;
			12'd1380: q <= 1'b0;
			12'd1381: q <= 1'b0;
			12'd1382: q <= 1'b0;
			12'd1383: q <= 1'b0;
			12'd1384: q <= 1'b0;
			12'd1385: q <= 1'b0;
			12'd1386: q <= 1'b0;
			12'd1387: q <= 1'b0;
			12'd1388: q <= 1'b1;
			12'd1389: q <= 1'b1;
			12'd1390: q <= 1'b1;
			12'd1391: q <= 1'b1;
			12'd1392: q <= 1'b1;
			12'd1393: q <= 1'b1;
			12'd1394: q <= 1'b1;
			12'd1395: q <= 1'b1;
			12'd1396: q <= 1'b1;
			12'd1397: q <= 1'b1;
			12'd1398: q <= 1'b1;
			12'd1399: q <= 1'b1;
			12'd1400: q <= 1'b1;
			12'd1401: q <= 1'b1;
			12'd1402: q <= 1'b1;
			12'd1403: q <= 1'b1;
			12'd1404: q <= 1'b1;
			12'd1405: q <= 1'b1;
			12'd1406: q <= 1'b1;
			12'd1407: q <= 1'b0;
			12'd1408: q <= 1'b0;
			12'd1409: q <= 1'b0;
			12'd1410: q <= 1'b0;
			12'd1411: q <= 1'b0;
			12'd1412: q <= 1'b0;
			12'd1413: q <= 1'b0;
			12'd1414: q <= 1'b0;
			12'd1415: q <= 1'b0;
			12'd1416: q <= 1'b0;
			12'd1417: q <= 1'b0;
			12'd1418: q <= 1'b0;
			12'd1419: q <= 1'b0;
			12'd1420: q <= 1'b0;
			12'd1421: q <= 1'b0;
			12'd1422: q <= 1'b0;
			12'd1423: q <= 1'b0;
			12'd1424: q <= 1'b0;
			12'd1425: q <= 1'b0;
			12'd1426: q <= 1'b0;
			12'd1427: q <= 1'b0;
			12'd1428: q <= 1'b1;
			12'd1429: q <= 1'b1;
			12'd1430: q <= 1'b1;
			12'd1431: q <= 1'b1;
			12'd1432: q <= 1'b1;
			12'd1433: q <= 1'b1;
			12'd1434: q <= 1'b1;
			12'd1435: q <= 1'b1;
			12'd1436: q <= 1'b1;
			12'd1437: q <= 1'b1;
			12'd1438: q <= 1'b1;
			12'd1439: q <= 1'b1;
			12'd1440: q <= 1'b1;
			12'd1441: q <= 1'b1;
			12'd1442: q <= 1'b1;
			12'd1443: q <= 1'b1;
			12'd1444: q <= 1'b1;
			12'd1445: q <= 1'b1;
			12'd1446: q <= 1'b1;
			12'd1447: q <= 1'b0;
			12'd1448: q <= 1'b0;
			12'd1449: q <= 1'b0;
			12'd1450: q <= 1'b0;
			12'd1451: q <= 1'b0;
			12'd1452: q <= 1'b0;
			12'd1453: q <= 1'b0;
			12'd1454: q <= 1'b0;
			12'd1455: q <= 1'b0;
			12'd1456: q <= 1'b0;
			12'd1457: q <= 1'b0;
			12'd1458: q <= 1'b0;
			12'd1459: q <= 1'b0;
			12'd1460: q <= 1'b0;
			12'd1461: q <= 1'b0;
			12'd1462: q <= 1'b0;
			12'd1463: q <= 1'b0;
			12'd1464: q <= 1'b0;
			12'd1465: q <= 1'b0;
			12'd1466: q <= 1'b0;
			12'd1467: q <= 1'b0;
			12'd1468: q <= 1'b1;
			12'd1469: q <= 1'b1;
			12'd1470: q <= 1'b1;
			12'd1471: q <= 1'b1;
			12'd1472: q <= 1'b1;
			12'd1473: q <= 1'b1;
			12'd1474: q <= 1'b1;
			12'd1475: q <= 1'b1;
			12'd1476: q <= 1'b1;
			12'd1477: q <= 1'b1;
			12'd1478: q <= 1'b1;
			12'd1479: q <= 1'b1;
			12'd1480: q <= 1'b1;
			12'd1481: q <= 1'b1;
			12'd1482: q <= 1'b1;
			12'd1483: q <= 1'b1;
			12'd1484: q <= 1'b1;
			12'd1485: q <= 1'b1;
			12'd1486: q <= 1'b1;
			12'd1487: q <= 1'b0;
			12'd1488: q <= 1'b0;
			12'd1489: q <= 1'b0;
			12'd1490: q <= 1'b0;
			12'd1491: q <= 1'b0;
			12'd1492: q <= 1'b0;
			12'd1493: q <= 1'b0;
			12'd1494: q <= 1'b0;
			12'd1495: q <= 1'b0;
			12'd1496: q <= 1'b0;
			12'd1497: q <= 1'b0;
			12'd1498: q <= 1'b0;
			12'd1499: q <= 1'b0;
			12'd1500: q <= 1'b0;
			12'd1501: q <= 1'b0;
			12'd1502: q <= 1'b0;
			12'd1503: q <= 1'b0;
			12'd1504: q <= 1'b0;
			12'd1505: q <= 1'b0;
			12'd1506: q <= 1'b0;
			12'd1507: q <= 1'b0;
			12'd1508: q <= 1'b1;
			12'd1509: q <= 1'b1;
			12'd1510: q <= 1'b1;
			12'd1511: q <= 1'b1;
			12'd1512: q <= 1'b1;
			12'd1513: q <= 1'b1;
			12'd1514: q <= 1'b1;
			12'd1515: q <= 1'b1;
			12'd1516: q <= 1'b1;
			12'd1517: q <= 1'b1;
			12'd1518: q <= 1'b1;
			12'd1519: q <= 1'b1;
			12'd1520: q <= 1'b1;
			12'd1521: q <= 1'b1;
			12'd1522: q <= 1'b1;
			12'd1523: q <= 1'b1;
			12'd1524: q <= 1'b1;
			12'd1525: q <= 1'b1;
			12'd1526: q <= 1'b1;
			12'd1527: q <= 1'b1;
			12'd1528: q <= 1'b0;
			12'd1529: q <= 1'b0;
			12'd1530: q <= 1'b0;
			12'd1531: q <= 1'b0;
			12'd1532: q <= 1'b0;
			12'd1533: q <= 1'b0;
			12'd1534: q <= 1'b0;
			12'd1535: q <= 1'b0;
			12'd1536: q <= 1'b0;
			12'd1537: q <= 1'b0;
			12'd1538: q <= 1'b0;
			12'd1539: q <= 1'b0;
			12'd1540: q <= 1'b0;
			12'd1541: q <= 1'b0;
			12'd1542: q <= 1'b0;
			12'd1543: q <= 1'b0;
			12'd1544: q <= 1'b0;
			12'd1545: q <= 1'b0;
			12'd1546: q <= 1'b0;
			12'd1547: q <= 1'b0;
			12'd1548: q <= 1'b1;
			12'd1549: q <= 1'b1;
			12'd1550: q <= 1'b1;
			12'd1551: q <= 1'b1;
			12'd1552: q <= 1'b1;
			12'd1553: q <= 1'b1;
			12'd1554: q <= 1'b1;
			12'd1555: q <= 1'b1;
			12'd1556: q <= 1'b1;
			12'd1557: q <= 1'b1;
			12'd1558: q <= 1'b1;
			12'd1559: q <= 1'b1;
			12'd1560: q <= 1'b1;
			12'd1561: q <= 1'b1;
			12'd1562: q <= 1'b1;
			12'd1563: q <= 1'b1;
			12'd1564: q <= 1'b1;
			12'd1565: q <= 1'b1;
			12'd1566: q <= 1'b1;
			12'd1567: q <= 1'b1;
			12'd1568: q <= 1'b0;
			12'd1569: q <= 1'b0;
			12'd1570: q <= 1'b0;
			12'd1571: q <= 1'b0;
			12'd1572: q <= 1'b0;
			12'd1573: q <= 1'b0;
			12'd1574: q <= 1'b0;
			12'd1575: q <= 1'b0;
			12'd1576: q <= 1'b0;
			12'd1577: q <= 1'b0;
			12'd1578: q <= 1'b0;
			12'd1579: q <= 1'b0;
			12'd1580: q <= 1'b0;
			12'd1581: q <= 1'b0;
			12'd1582: q <= 1'b0;
			12'd1583: q <= 1'b0;
			12'd1584: q <= 1'b0;
			12'd1585: q <= 1'b0;
			12'd1586: q <= 1'b0;
			12'd1587: q <= 1'b0;
			12'd1588: q <= 1'b1;
			12'd1589: q <= 1'b1;
			12'd1590: q <= 1'b1;
			12'd1591: q <= 1'b1;
			12'd1592: q <= 1'b1;
			12'd1593: q <= 1'b1;
			12'd1594: q <= 1'b1;
			12'd1595: q <= 1'b1;
			12'd1596: q <= 1'b1;
			12'd1597: q <= 1'b1;
			12'd1598: q <= 1'b1;
			12'd1599: q <= 1'b1;
			12'd1600: q <= 1'b1;
			12'd1601: q <= 1'b1;
			12'd1602: q <= 1'b1;
			12'd1603: q <= 1'b1;
			12'd1604: q <= 1'b1;
			12'd1605: q <= 1'b1;
			12'd1606: q <= 1'b1;
			12'd1607: q <= 1'b1;
			12'd1608: q <= 1'b0;
			12'd1609: q <= 1'b0;
			12'd1610: q <= 1'b0;
			12'd1611: q <= 1'b0;
			12'd1612: q <= 1'b0;
			12'd1613: q <= 1'b0;
			12'd1614: q <= 1'b0;
			12'd1615: q <= 1'b0;
			12'd1616: q <= 1'b0;
			12'd1617: q <= 1'b0;
			12'd1618: q <= 1'b0;
			12'd1619: q <= 1'b0;
			12'd1620: q <= 1'b0;
			12'd1621: q <= 1'b0;
			12'd1622: q <= 1'b0;
			12'd1623: q <= 1'b0;
			12'd1624: q <= 1'b0;
			12'd1625: q <= 1'b0;
			12'd1626: q <= 1'b0;
			12'd1627: q <= 1'b1;
			12'd1628: q <= 1'b1;
			12'd1629: q <= 1'b1;
			12'd1630: q <= 1'b1;
			12'd1631: q <= 1'b1;
			12'd1632: q <= 1'b1;
			12'd1633: q <= 1'b1;
			12'd1634: q <= 1'b1;
			12'd1635: q <= 1'b1;
			12'd1636: q <= 1'b1;
			12'd1637: q <= 1'b1;
			12'd1638: q <= 1'b1;
			12'd1639: q <= 1'b1;
			12'd1640: q <= 1'b1;
			12'd1641: q <= 1'b1;
			12'd1642: q <= 1'b1;
			12'd1643: q <= 1'b1;
			12'd1644: q <= 1'b1;
			12'd1645: q <= 1'b1;
			12'd1646: q <= 1'b1;
			12'd1647: q <= 1'b1;
			12'd1648: q <= 1'b0;
			12'd1649: q <= 1'b0;
			12'd1650: q <= 1'b0;
			12'd1651: q <= 1'b0;
			12'd1652: q <= 1'b0;
			12'd1653: q <= 1'b0;
			12'd1654: q <= 1'b0;
			12'd1655: q <= 1'b0;
			12'd1656: q <= 1'b0;
			12'd1657: q <= 1'b0;
			12'd1658: q <= 1'b0;
			12'd1659: q <= 1'b0;
			12'd1660: q <= 1'b0;
			12'd1661: q <= 1'b0;
			12'd1662: q <= 1'b0;
			12'd1663: q <= 1'b0;
			12'd1664: q <= 1'b0;
			12'd1665: q <= 1'b0;
			12'd1666: q <= 1'b0;
			12'd1667: q <= 1'b1;
			12'd1668: q <= 1'b1;
			12'd1669: q <= 1'b1;
			12'd1670: q <= 1'b1;
			12'd1671: q <= 1'b1;
			12'd1672: q <= 1'b1;
			12'd1673: q <= 1'b1;
			12'd1674: q <= 1'b1;
			12'd1675: q <= 1'b1;
			12'd1676: q <= 1'b1;
			12'd1677: q <= 1'b1;
			12'd1678: q <= 1'b1;
			12'd1679: q <= 1'b1;
			12'd1680: q <= 1'b1;
			12'd1681: q <= 1'b1;
			12'd1682: q <= 1'b1;
			12'd1683: q <= 1'b1;
			12'd1684: q <= 1'b1;
			12'd1685: q <= 1'b1;
			12'd1686: q <= 1'b1;
			12'd1687: q <= 1'b1;
			12'd1688: q <= 1'b1;
			12'd1689: q <= 1'b0;
			12'd1690: q <= 1'b0;
			12'd1691: q <= 1'b0;
			12'd1692: q <= 1'b0;
			12'd1693: q <= 1'b0;
			12'd1694: q <= 1'b0;
			12'd1695: q <= 1'b0;
			12'd1696: q <= 1'b0;
			12'd1697: q <= 1'b0;
			12'd1698: q <= 1'b0;
			12'd1699: q <= 1'b0;
			12'd1700: q <= 1'b0;
			12'd1701: q <= 1'b0;
			12'd1702: q <= 1'b0;
			12'd1703: q <= 1'b0;
			12'd1704: q <= 1'b0;
			12'd1705: q <= 1'b0;
			12'd1706: q <= 1'b0;
			12'd1707: q <= 1'b0;
			12'd1708: q <= 1'b1;
			12'd1709: q <= 1'b1;
			12'd1710: q <= 1'b1;
			12'd1711: q <= 1'b1;
			12'd1712: q <= 1'b1;
			12'd1713: q <= 1'b1;
			12'd1714: q <= 1'b1;
			12'd1715: q <= 1'b1;
			12'd1716: q <= 1'b1;
			12'd1717: q <= 1'b1;
			12'd1718: q <= 1'b1;
			12'd1719: q <= 1'b1;
			12'd1720: q <= 1'b1;
			12'd1721: q <= 1'b1;
			12'd1722: q <= 1'b1;
			12'd1723: q <= 1'b1;
			12'd1724: q <= 1'b1;
			12'd1725: q <= 1'b1;
			12'd1726: q <= 1'b1;
			12'd1727: q <= 1'b1;
			12'd1728: q <= 1'b1;
			12'd1729: q <= 1'b0;
			12'd1730: q <= 1'b0;
			12'd1731: q <= 1'b0;
			12'd1732: q <= 1'b0;
			12'd1733: q <= 1'b0;
			12'd1734: q <= 1'b0;
			12'd1735: q <= 1'b0;
			12'd1736: q <= 1'b0;
			12'd1737: q <= 1'b0;
			12'd1738: q <= 1'b0;
			12'd1739: q <= 1'b0;
			12'd1740: q <= 1'b0;
			12'd1741: q <= 1'b0;
			12'd1742: q <= 1'b0;
			12'd1743: q <= 1'b0;
			12'd1744: q <= 1'b0;
			12'd1745: q <= 1'b0;
			12'd1746: q <= 1'b0;
			12'd1747: q <= 1'b0;
			12'd1748: q <= 1'b1;
			12'd1749: q <= 1'b1;
			12'd1750: q <= 1'b1;
			12'd1751: q <= 1'b1;
			12'd1752: q <= 1'b1;
			12'd1753: q <= 1'b1;
			12'd1754: q <= 1'b1;
			12'd1755: q <= 1'b1;
			12'd1756: q <= 1'b1;
			12'd1757: q <= 1'b1;
			12'd1758: q <= 1'b1;
			12'd1759: q <= 1'b1;
			12'd1760: q <= 1'b1;
			12'd1761: q <= 1'b1;
			12'd1762: q <= 1'b1;
			12'd1763: q <= 1'b1;
			12'd1764: q <= 1'b1;
			12'd1765: q <= 1'b1;
			12'd1766: q <= 1'b1;
			12'd1767: q <= 1'b1;
			12'd1768: q <= 1'b1;
			12'd1769: q <= 1'b1;
			12'd1770: q <= 1'b0;
			12'd1771: q <= 1'b0;
			12'd1772: q <= 1'b0;
			12'd1773: q <= 1'b0;
			12'd1774: q <= 1'b0;
			12'd1775: q <= 1'b0;
			12'd1776: q <= 1'b0;
			12'd1777: q <= 1'b0;
			12'd1778: q <= 1'b0;
			12'd1779: q <= 1'b0;
			12'd1780: q <= 1'b0;
			12'd1781: q <= 1'b0;
			12'd1782: q <= 1'b0;
			12'd1783: q <= 1'b0;
			12'd1784: q <= 1'b0;
			12'd1785: q <= 1'b0;
			12'd1786: q <= 1'b0;
			12'd1787: q <= 1'b0;
			12'd1788: q <= 1'b0;
			12'd1789: q <= 1'b0;
			12'd1790: q <= 1'b0;
			12'd1791: q <= 1'b0;
			12'd1792: q <= 1'b1;
			12'd1793: q <= 1'b1;
			12'd1794: q <= 1'b1;
			12'd1795: q <= 1'b1;
			12'd1796: q <= 1'b1;
			12'd1797: q <= 1'b1;
			12'd1798: q <= 1'b1;
			12'd1799: q <= 1'b1;
			12'd1800: q <= 1'b1;
			12'd1801: q <= 1'b1;
			12'd1802: q <= 1'b1;
			12'd1803: q <= 1'b1;
			12'd1804: q <= 1'b1;
			12'd1805: q <= 1'b1;
			12'd1806: q <= 1'b1;
			12'd1807: q <= 1'b1;
			12'd1808: q <= 1'b1;
			12'd1809: q <= 1'b1;
			12'd1810: q <= 1'b0;
			12'd1811: q <= 1'b0;
			12'd1812: q <= 1'b0;
			12'd1813: q <= 1'b0;
			12'd1814: q <= 1'b0;
			12'd1815: q <= 1'b0;
			12'd1816: q <= 1'b0;
			12'd1817: q <= 1'b0;
			12'd1818: q <= 1'b0;
			12'd1819: q <= 1'b0;
			12'd1820: q <= 1'b0;
			12'd1821: q <= 1'b0;
			12'd1822: q <= 1'b0;
			12'd1823: q <= 1'b0;
			12'd1824: q <= 1'b0;
			12'd1825: q <= 1'b0;
			12'd1826: q <= 1'b0;
			12'd1827: q <= 1'b0;
			12'd1828: q <= 1'b0;
			12'd1829: q <= 1'b0;
			12'd1830: q <= 1'b0;
			12'd1831: q <= 1'b0;
			12'd1832: q <= 1'b0;
			12'd1833: q <= 1'b0;
			12'd1834: q <= 1'b1;
			12'd1835: q <= 1'b1;
			12'd1836: q <= 1'b1;
			12'd1837: q <= 1'b1;
			12'd1838: q <= 1'b1;
			12'd1839: q <= 1'b1;
			12'd1840: q <= 1'b1;
			12'd1841: q <= 1'b1;
			12'd1842: q <= 1'b1;
			12'd1843: q <= 1'b1;
			12'd1844: q <= 1'b1;
			12'd1845: q <= 1'b1;
			12'd1846: q <= 1'b1;
			12'd1847: q <= 1'b1;
			12'd1848: q <= 1'b1;
			12'd1849: q <= 1'b1;
			12'd1850: q <= 1'b0;
			12'd1851: q <= 1'b0;
			12'd1852: q <= 1'b0;
			12'd1853: q <= 1'b0;
			12'd1854: q <= 1'b0;
			12'd1855: q <= 1'b0;
			12'd1856: q <= 1'b0;
			12'd1857: q <= 1'b0;
			12'd1858: q <= 1'b0;
			12'd1859: q <= 1'b0;
			12'd1860: q <= 1'b0;
			12'd1861: q <= 1'b0;
			12'd1862: q <= 1'b0;
			12'd1863: q <= 1'b0;
			12'd1864: q <= 1'b0;
			12'd1865: q <= 1'b0;
			12'd1866: q <= 1'b0;
			12'd1867: q <= 1'b0;
			12'd1868: q <= 1'b0;
			12'd1869: q <= 1'b0;
			12'd1870: q <= 1'b0;
			12'd1871: q <= 1'b0;
			12'd1872: q <= 1'b0;
			12'd1873: q <= 1'b0;
			12'd1874: q <= 1'b0;
			12'd1875: q <= 1'b0;
			12'd1876: q <= 1'b0;
			12'd1877: q <= 1'b0;
			12'd1878: q <= 1'b0;
			12'd1879: q <= 1'b0;
			12'd1880: q <= 1'b1;
			12'd1881: q <= 1'b1;
			12'd1882: q <= 1'b1;
			12'd1883: q <= 1'b1;
			12'd1884: q <= 1'b1;
			12'd1885: q <= 1'b1;
			12'd1886: q <= 1'b1;
			12'd1887: q <= 1'b1;
			12'd1888: q <= 1'b1;
			12'd1889: q <= 1'b1;
			12'd1890: q <= 1'b0;
			12'd1891: q <= 1'b0;
			12'd1892: q <= 1'b0;
			12'd1893: q <= 1'b0;
			12'd1894: q <= 1'b0;
			12'd1895: q <= 1'b0;
			12'd1896: q <= 1'b0;
			12'd1897: q <= 1'b0;
			12'd1898: q <= 1'b0;
			12'd1899: q <= 1'b0;
			12'd1900: q <= 1'b0;
			12'd1901: q <= 1'b0;
			12'd1902: q <= 1'b0;
			12'd1903: q <= 1'b0;
			12'd1904: q <= 1'b0;
			12'd1905: q <= 1'b0;
			12'd1906: q <= 1'b0;
			12'd1907: q <= 1'b0;
			12'd1908: q <= 1'b0;
			12'd1909: q <= 1'b1;
			12'd1910: q <= 1'b0;
			12'd1911: q <= 1'b0;
			12'd1912: q <= 1'b0;
			12'd1913: q <= 1'b0;
			12'd1914: q <= 1'b0;
			12'd1915: q <= 1'b0;
			12'd1916: q <= 1'b1;
			12'd1917: q <= 1'b1;
			12'd1918: q <= 1'b1;
			12'd1919: q <= 1'b1;
			12'd1920: q <= 1'b1;
			12'd1921: q <= 1'b1;
			12'd1922: q <= 1'b1;
			12'd1923: q <= 1'b1;
			12'd1924: q <= 1'b1;
			12'd1925: q <= 1'b1;
			12'd1926: q <= 1'b1;
			12'd1927: q <= 1'b1;
			12'd1928: q <= 1'b1;
			12'd1929: q <= 1'b0;
			12'd1930: q <= 1'b0;
			12'd1931: q <= 1'b0;
			12'd1932: q <= 1'b0;
			12'd1933: q <= 1'b0;
			12'd1934: q <= 1'b0;
			12'd1935: q <= 1'b0;
			12'd1936: q <= 1'b0;
			12'd1937: q <= 1'b0;
			12'd1938: q <= 1'b0;
			12'd1939: q <= 1'b0;
			12'd1940: q <= 1'b0;
			12'd1941: q <= 1'b0;
			12'd1942: q <= 1'b0;
			12'd1943: q <= 1'b0;
			12'd1944: q <= 1'b0;
			12'd1945: q <= 1'b0;
			12'd1946: q <= 1'b0;
			12'd1947: q <= 1'b0;
			12'd1948: q <= 1'b0;
			12'd1949: q <= 1'b1;
			12'd1950: q <= 1'b1;
			12'd1951: q <= 1'b1;
			12'd1952: q <= 1'b0;
			12'd1953: q <= 1'b0;
			12'd1954: q <= 1'b1;
			12'd1955: q <= 1'b1;
			12'd1956: q <= 1'b1;
			12'd1957: q <= 1'b1;
			12'd1958: q <= 1'b1;
			12'd1959: q <= 1'b1;
			12'd1960: q <= 1'b1;
			12'd1961: q <= 1'b1;
			12'd1962: q <= 1'b1;
			12'd1963: q <= 1'b1;
			12'd1964: q <= 1'b1;
			12'd1965: q <= 1'b1;
			12'd1966: q <= 1'b1;
			12'd1967: q <= 1'b1;
			12'd1968: q <= 1'b1;
			12'd1969: q <= 1'b1;
			12'd1970: q <= 1'b0;
			12'd1971: q <= 1'b0;
			12'd1972: q <= 1'b0;
			12'd1973: q <= 1'b0;
			12'd1974: q <= 1'b0;
			12'd1975: q <= 1'b0;
			12'd1976: q <= 1'b0;
			12'd1977: q <= 1'b0;
			12'd1978: q <= 1'b0;
			12'd1979: q <= 1'b0;
			12'd1980: q <= 1'b0;
			12'd1981: q <= 1'b0;
			12'd1982: q <= 1'b0;
			12'd1983: q <= 1'b0;
			12'd1984: q <= 1'b0;
			12'd1985: q <= 1'b0;
			12'd1986: q <= 1'b0;
			12'd1987: q <= 1'b0;
			12'd1988: q <= 1'b0;
			12'd1989: q <= 1'b0;
			12'd1990: q <= 1'b1;
			12'd1991: q <= 1'b1;
			12'd1992: q <= 1'b1;
			12'd1993: q <= 1'b1;
			12'd1994: q <= 1'b1;
			12'd1995: q <= 1'b1;
			12'd1996: q <= 1'b1;
			12'd1997: q <= 1'b1;
			12'd1998: q <= 1'b1;
			12'd1999: q <= 1'b1;
			12'd2000: q <= 1'b1;
			12'd2001: q <= 1'b1;
			12'd2002: q <= 1'b1;
			12'd2003: q <= 1'b1;
			12'd2004: q <= 1'b1;
			12'd2005: q <= 1'b1;
			12'd2006: q <= 1'b1;
			12'd2007: q <= 1'b1;
			12'd2008: q <= 1'b1;
			12'd2009: q <= 1'b1;
			12'd2010: q <= 1'b0;
			12'd2011: q <= 1'b0;
			12'd2012: q <= 1'b0;
			12'd2013: q <= 1'b0;
			12'd2014: q <= 1'b0;
			12'd2015: q <= 1'b0;
			12'd2016: q <= 1'b0;
			12'd2017: q <= 1'b0;
			12'd2018: q <= 1'b0;
			12'd2019: q <= 1'b0;
			12'd2020: q <= 1'b0;
			12'd2021: q <= 1'b0;
			12'd2022: q <= 1'b0;
			12'd2023: q <= 1'b0;
			12'd2024: q <= 1'b0;
			12'd2025: q <= 1'b0;
			12'd2026: q <= 1'b0;
			12'd2027: q <= 1'b0;
			12'd2028: q <= 1'b0;
			12'd2029: q <= 1'b0;
			12'd2030: q <= 1'b0;
			12'd2031: q <= 1'b1;
			12'd2032: q <= 1'b1;
			12'd2033: q <= 1'b1;
			12'd2034: q <= 1'b1;
			12'd2035: q <= 1'b1;
			12'd2036: q <= 1'b1;
			12'd2037: q <= 1'b1;
			12'd2038: q <= 1'b1;
			12'd2039: q <= 1'b1;
			12'd2040: q <= 1'b1;
			12'd2041: q <= 1'b1;
			12'd2042: q <= 1'b1;
			12'd2043: q <= 1'b1;
			12'd2044: q <= 1'b1;
			12'd2045: q <= 1'b1;
			12'd2046: q <= 1'b1;
			12'd2047: q <= 1'b1;
			12'd2048: q <= 1'b1;
			12'd2049: q <= 1'b1;
			12'd2050: q <= 1'b0;
			12'd2051: q <= 1'b0;
			12'd2052: q <= 1'b0;
			12'd2053: q <= 1'b0;
			12'd2054: q <= 1'b0;
			12'd2055: q <= 1'b0;
			12'd2056: q <= 1'b0;
			12'd2057: q <= 1'b0;
			12'd2058: q <= 1'b0;
			12'd2059: q <= 1'b0;
			12'd2060: q <= 1'b0;
			12'd2061: q <= 1'b0;
			12'd2062: q <= 1'b0;
			12'd2063: q <= 1'b0;
			12'd2064: q <= 1'b0;
			12'd2065: q <= 1'b0;
			12'd2066: q <= 1'b0;
			12'd2067: q <= 1'b0;
			12'd2068: q <= 1'b0;
			12'd2069: q <= 1'b0;
			12'd2070: q <= 1'b1;
			12'd2071: q <= 1'b1;
			12'd2072: q <= 1'b1;
			12'd2073: q <= 1'b1;
			12'd2074: q <= 1'b1;
			12'd2075: q <= 1'b1;
			12'd2076: q <= 1'b1;
			12'd2077: q <= 1'b1;
			12'd2078: q <= 1'b1;
			12'd2079: q <= 1'b1;
			12'd2080: q <= 1'b1;
			12'd2081: q <= 1'b1;
			12'd2082: q <= 1'b1;
			12'd2083: q <= 1'b1;
			12'd2084: q <= 1'b1;
			12'd2085: q <= 1'b1;
			12'd2086: q <= 1'b1;
			12'd2087: q <= 1'b1;
			12'd2088: q <= 1'b1;
			12'd2089: q <= 1'b0;
			12'd2090: q <= 1'b0;
			12'd2091: q <= 1'b0;
			12'd2092: q <= 1'b0;
			12'd2093: q <= 1'b0;
			12'd2094: q <= 1'b0;
			12'd2095: q <= 1'b0;
			12'd2096: q <= 1'b0;
			12'd2097: q <= 1'b0;
			12'd2098: q <= 1'b0;
			12'd2099: q <= 1'b0;
			12'd2100: q <= 1'b0;
			12'd2101: q <= 1'b0;
			12'd2102: q <= 1'b0;
			12'd2103: q <= 1'b0;
			12'd2104: q <= 1'b0;
			12'd2105: q <= 1'b0;
			12'd2106: q <= 1'b0;
			12'd2107: q <= 1'b0;
			12'd2108: q <= 1'b0;
			12'd2109: q <= 1'b0;
			12'd2110: q <= 1'b0;
			12'd2111: q <= 1'b1;
			12'd2112: q <= 1'b1;
			12'd2113: q <= 1'b1;
			12'd2114: q <= 1'b1;
			12'd2115: q <= 1'b1;
			12'd2116: q <= 1'b1;
			12'd2117: q <= 1'b1;
			12'd2118: q <= 1'b1;
			12'd2119: q <= 1'b1;
			12'd2120: q <= 1'b1;
			12'd2121: q <= 1'b1;
			12'd2122: q <= 1'b1;
			12'd2123: q <= 1'b1;
			12'd2124: q <= 1'b1;
			12'd2125: q <= 1'b1;
			12'd2126: q <= 1'b1;
			12'd2127: q <= 1'b1;
			12'd2128: q <= 1'b1;
			12'd2129: q <= 1'b0;
			12'd2130: q <= 1'b0;
			12'd2131: q <= 1'b0;
			12'd2132: q <= 1'b0;
			12'd2133: q <= 1'b0;
			12'd2134: q <= 1'b0;
			12'd2135: q <= 1'b0;
			12'd2136: q <= 1'b0;
			12'd2137: q <= 1'b0;
			12'd2138: q <= 1'b0;
			12'd2139: q <= 1'b0;
			12'd2140: q <= 1'b0;
			12'd2141: q <= 1'b0;
			12'd2142: q <= 1'b0;
			12'd2143: q <= 1'b0;
			12'd2144: q <= 1'b0;
			12'd2145: q <= 1'b0;
			12'd2146: q <= 1'b0;
			12'd2147: q <= 1'b0;
			12'd2148: q <= 1'b0;
			12'd2149: q <= 1'b0;
			12'd2150: q <= 1'b0;
			12'd2151: q <= 1'b1;
			12'd2152: q <= 1'b1;
			12'd2153: q <= 1'b1;
			12'd2154: q <= 1'b1;
			12'd2155: q <= 1'b1;
			12'd2156: q <= 1'b1;
			12'd2157: q <= 1'b1;
			12'd2158: q <= 1'b1;
			12'd2159: q <= 1'b1;
			12'd2160: q <= 1'b1;
			12'd2161: q <= 1'b1;
			12'd2162: q <= 1'b1;
			12'd2163: q <= 1'b1;
			12'd2164: q <= 1'b1;
			12'd2165: q <= 1'b1;
			12'd2166: q <= 1'b1;
			12'd2167: q <= 1'b1;
			12'd2168: q <= 1'b1;
			12'd2169: q <= 1'b0;
			12'd2170: q <= 1'b0;
			12'd2171: q <= 1'b0;
			12'd2172: q <= 1'b0;
			12'd2173: q <= 1'b0;
			12'd2174: q <= 1'b0;
			12'd2175: q <= 1'b0;
			12'd2176: q <= 1'b0;
			12'd2177: q <= 1'b0;
			12'd2178: q <= 1'b0;
			12'd2179: q <= 1'b0;
			12'd2180: q <= 1'b0;
			12'd2181: q <= 1'b0;
			12'd2182: q <= 1'b0;
			12'd2183: q <= 1'b0;
			12'd2184: q <= 1'b0;
			12'd2185: q <= 1'b0;
			12'd2186: q <= 1'b0;
			12'd2187: q <= 1'b0;
			12'd2188: q <= 1'b0;
			12'd2189: q <= 1'b0;
			12'd2190: q <= 1'b0;
			12'd2191: q <= 1'b1;
			12'd2192: q <= 1'b1;
			12'd2193: q <= 1'b1;
			12'd2194: q <= 1'b1;
			12'd2195: q <= 1'b1;
			12'd2196: q <= 1'b1;
			12'd2197: q <= 1'b1;
			12'd2198: q <= 1'b1;
			12'd2199: q <= 1'b1;
			12'd2200: q <= 1'b1;
			12'd2201: q <= 1'b1;
			12'd2202: q <= 1'b1;
			12'd2203: q <= 1'b1;
			12'd2204: q <= 1'b1;
			12'd2205: q <= 1'b1;
			12'd2206: q <= 1'b1;
			12'd2207: q <= 1'b1;
			12'd2208: q <= 1'b1;
			12'd2209: q <= 1'b0;
			12'd2210: q <= 1'b0;
			12'd2211: q <= 1'b0;
			12'd2212: q <= 1'b0;
			12'd2213: q <= 1'b0;
			12'd2214: q <= 1'b0;
			12'd2215: q <= 1'b0;
			12'd2216: q <= 1'b0;
			12'd2217: q <= 1'b0;
			12'd2218: q <= 1'b0;
			12'd2219: q <= 1'b0;
			12'd2220: q <= 1'b0;
			12'd2221: q <= 1'b0;
			12'd2222: q <= 1'b0;
			12'd2223: q <= 1'b0;
			12'd2224: q <= 1'b0;
			12'd2225: q <= 1'b0;
			12'd2226: q <= 1'b0;
			12'd2227: q <= 1'b0;
			12'd2228: q <= 1'b0;
			12'd2229: q <= 1'b0;
			12'd2230: q <= 1'b0;
			12'd2231: q <= 1'b1;
			12'd2232: q <= 1'b1;
			12'd2233: q <= 1'b1;
			12'd2234: q <= 1'b1;
			12'd2235: q <= 1'b1;
			12'd2236: q <= 1'b1;
			12'd2237: q <= 1'b1;
			12'd2238: q <= 1'b1;
			12'd2239: q <= 1'b1;
			12'd2240: q <= 1'b1;
			12'd2241: q <= 1'b1;
			12'd2242: q <= 1'b1;
			12'd2243: q <= 1'b1;
			12'd2244: q <= 1'b1;
			12'd2245: q <= 1'b1;
			12'd2246: q <= 1'b1;
			12'd2247: q <= 1'b1;
			12'd2248: q <= 1'b1;
			12'd2249: q <= 1'b0;
			12'd2250: q <= 1'b0;
			12'd2251: q <= 1'b0;
			12'd2252: q <= 1'b0;
			12'd2253: q <= 1'b0;
			12'd2254: q <= 1'b0;
			12'd2255: q <= 1'b0;
			12'd2256: q <= 1'b0;
			12'd2257: q <= 1'b0;
			12'd2258: q <= 1'b0;
			12'd2259: q <= 1'b0;
			12'd2260: q <= 1'b0;
			12'd2261: q <= 1'b0;
			12'd2262: q <= 1'b0;
			12'd2263: q <= 1'b0;
			12'd2264: q <= 1'b0;
			12'd2265: q <= 1'b0;
			12'd2266: q <= 1'b0;
			12'd2267: q <= 1'b0;
			12'd2268: q <= 1'b0;
			12'd2269: q <= 1'b0;
			12'd2270: q <= 1'b0;
			12'd2271: q <= 1'b1;
			12'd2272: q <= 1'b1;
			12'd2273: q <= 1'b1;
			12'd2274: q <= 1'b1;
			12'd2275: q <= 1'b1;
			12'd2276: q <= 1'b1;
			12'd2277: q <= 1'b1;
			12'd2278: q <= 1'b1;
			12'd2279: q <= 1'b1;
			12'd2280: q <= 1'b1;
			12'd2281: q <= 1'b1;
			12'd2282: q <= 1'b1;
			12'd2283: q <= 1'b1;
			12'd2284: q <= 1'b1;
			12'd2285: q <= 1'b1;
			12'd2286: q <= 1'b1;
			12'd2287: q <= 1'b1;
			12'd2288: q <= 1'b1;
			12'd2289: q <= 1'b1;
			12'd2290: q <= 1'b0;
			12'd2291: q <= 1'b0;
			12'd2292: q <= 1'b0;
			12'd2293: q <= 1'b0;
			12'd2294: q <= 1'b0;
			12'd2295: q <= 1'b0;
			12'd2296: q <= 1'b0;
			12'd2297: q <= 1'b0;
			12'd2298: q <= 1'b0;
			12'd2299: q <= 1'b0;
			12'd2300: q <= 1'b0;
			12'd2301: q <= 1'b0;
			12'd2302: q <= 1'b0;
			12'd2303: q <= 1'b0;
			12'd2304: q <= 1'b0;
			12'd2305: q <= 1'b0;
			12'd2306: q <= 1'b0;
			12'd2307: q <= 1'b0;
			12'd2308: q <= 1'b0;
			12'd2309: q <= 1'b0;
			12'd2310: q <= 1'b0;
			12'd2311: q <= 1'b1;
			12'd2312: q <= 1'b1;
			12'd2313: q <= 1'b1;
			12'd2314: q <= 1'b1;
			12'd2315: q <= 1'b1;
			12'd2316: q <= 1'b1;
			12'd2317: q <= 1'b1;
			12'd2318: q <= 1'b1;
			12'd2319: q <= 1'b1;
			12'd2320: q <= 1'b0;
			12'd2321: q <= 1'b0;
			12'd2322: q <= 1'b0;
			12'd2323: q <= 1'b0;
			12'd2324: q <= 1'b0;
			12'd2325: q <= 1'b0;
			12'd2326: q <= 1'b0;
			12'd2327: q <= 1'b0;
			12'd2328: q <= 1'b0;
			12'd2329: q <= 1'b0;
			12'd2330: q <= 1'b0;
			12'd2331: q <= 1'b0;
			12'd2332: q <= 1'b0;
			12'd2333: q <= 1'b0;
			12'd2334: q <= 1'b0;
			12'd2335: q <= 1'b0;
			12'd2336: q <= 1'b0;
			12'd2337: q <= 1'b0;
			12'd2338: q <= 1'b0;
			12'd2339: q <= 1'b0;
			12'd2340: q <= 1'b0;
			12'd2341: q <= 1'b0;
			12'd2342: q <= 1'b0;
			12'd2343: q <= 1'b0;
			12'd2344: q <= 1'b0;
			12'd2345: q <= 1'b0;
			12'd2346: q <= 1'b0;
			12'd2347: q <= 1'b0;
			12'd2348: q <= 1'b0;
			12'd2349: q <= 1'b0;
			12'd2350: q <= 1'b0;
			12'd2351: q <= 1'b0;
			12'd2352: q <= 1'b1;
			12'd2353: q <= 1'b1;
			12'd2354: q <= 1'b1;
			12'd2355: q <= 1'b1;
			12'd2356: q <= 1'b1;
			12'd2357: q <= 1'b1;
			12'd2358: q <= 1'b1;
			12'd2359: q <= 1'b1;
			12'd2360: q <= 1'b0;
			12'd2361: q <= 1'b0;
			12'd2362: q <= 1'b0;
			12'd2363: q <= 1'b0;
			12'd2364: q <= 1'b0;
			12'd2365: q <= 1'b0;
			12'd2366: q <= 1'b0;
			12'd2367: q <= 1'b0;
			12'd2368: q <= 1'b0;
			12'd2369: q <= 1'b0;
			12'd2370: q <= 1'b0;
			12'd2371: q <= 1'b0;
			12'd2372: q <= 1'b0;
			12'd2373: q <= 1'b0;
			12'd2374: q <= 1'b0;
			12'd2375: q <= 1'b0;
			12'd2376: q <= 1'b0;
			12'd2377: q <= 1'b0;
			12'd2378: q <= 1'b0;
			12'd2379: q <= 1'b0;
			12'd2380: q <= 1'b0;
			12'd2381: q <= 1'b0;
			12'd2382: q <= 1'b0;
			12'd2383: q <= 1'b0;
			12'd2384: q <= 1'b0;
			12'd2385: q <= 1'b0;
			12'd2386: q <= 1'b0;
			12'd2387: q <= 1'b0;
			12'd2388: q <= 1'b0;
			12'd2389: q <= 1'b0;
			12'd2390: q <= 1'b0;
			12'd2391: q <= 1'b0;
			12'd2392: q <= 1'b0;
			12'd2393: q <= 1'b0;
			12'd2394: q <= 1'b0;
			12'd2395: q <= 1'b0;
			12'd2396: q <= 1'b0;
			12'd2397: q <= 1'b0;
			12'd2398: q <= 1'b0;
			12'd2399: q <= 1'b0;
			12'd2400: q <= 1'b0;
			12'd2401: q <= 1'b0;
			12'd2402: q <= 1'b0;
			12'd2403: q <= 1'b0;
			12'd2404: q <= 1'b0;
			12'd2405: q <= 1'b0;
			12'd2406: q <= 1'b0;
			12'd2407: q <= 1'b0;
			12'd2408: q <= 1'b0;
			12'd2409: q <= 1'b0;
			12'd2410: q <= 1'b0;
			12'd2411: q <= 1'b0;
			12'd2412: q <= 1'b0;
			12'd2413: q <= 1'b0;
			12'd2414: q <= 1'b0;
			12'd2415: q <= 1'b0;
			12'd2416: q <= 1'b0;
			12'd2417: q <= 1'b0;
			12'd2418: q <= 1'b0;
			12'd2419: q <= 1'b0;
			12'd2420: q <= 1'b0;
			12'd2421: q <= 1'b0;
			12'd2422: q <= 1'b0;
			12'd2423: q <= 1'b0;
			12'd2424: q <= 1'b0;
			12'd2425: q <= 1'b0;
			12'd2426: q <= 1'b0;
			12'd2427: q <= 1'b0;
			12'd2428: q <= 1'b0;
			12'd2429: q <= 1'b0;
			12'd2430: q <= 1'b0;
			12'd2431: q <= 1'b0;
			12'd2432: q <= 1'b0;
			12'd2433: q <= 1'b0;
			12'd2434: q <= 1'b0;
			12'd2435: q <= 1'b0;
			12'd2436: q <= 1'b0;
			12'd2437: q <= 1'b0;
			12'd2438: q <= 1'b0;
			12'd2439: q <= 1'b0;
			12'd2440: q <= 1'b0;
			12'd2441: q <= 1'b0;
			12'd2442: q <= 1'b0;
			12'd2443: q <= 1'b0;
			12'd2444: q <= 1'b0;
			12'd2445: q <= 1'b0;
			12'd2446: q <= 1'b0;
			12'd2447: q <= 1'b0;
			12'd2448: q <= 1'b0;
			12'd2449: q <= 1'b0;
			12'd2450: q <= 1'b0;
			12'd2451: q <= 1'b0;
			12'd2452: q <= 1'b0;
			12'd2453: q <= 1'b0;
			12'd2454: q <= 1'b0;
			12'd2455: q <= 1'b0;
			12'd2456: q <= 1'b0;
			12'd2457: q <= 1'b0;
			12'd2458: q <= 1'b0;
			12'd2459: q <= 1'b0;
			12'd2460: q <= 1'b0;
			12'd2461: q <= 1'b0;
			12'd2462: q <= 1'b0;
			12'd2463: q <= 1'b0;
			12'd2464: q <= 1'b0;
			12'd2465: q <= 1'b0;
			12'd2466: q <= 1'b0;
			12'd2467: q <= 1'b0;
			12'd2468: q <= 1'b0;
			12'd2469: q <= 1'b0;
			12'd2470: q <= 1'b0;
			12'd2471: q <= 1'b0;
			12'd2472: q <= 1'b0;
			12'd2473: q <= 1'b0;
			12'd2474: q <= 1'b0;
			12'd2475: q <= 1'b0;
			12'd2476: q <= 1'b0;
			12'd2477: q <= 1'b0;
			12'd2478: q <= 1'b0;
			12'd2479: q <= 1'b0;
			12'd2480: q <= 1'b0;
			12'd2481: q <= 1'b0;
			12'd2482: q <= 1'b0;
			12'd2483: q <= 1'b0;
			12'd2484: q <= 1'b0;
			12'd2485: q <= 1'b0;
			12'd2486: q <= 1'b0;
			12'd2487: q <= 1'b0;
			12'd2488: q <= 1'b0;
			12'd2489: q <= 1'b0;
			12'd2490: q <= 1'b0;
			12'd2491: q <= 1'b0;
			12'd2492: q <= 1'b0;
			12'd2493: q <= 1'b0;
			12'd2494: q <= 1'b0;
			12'd2495: q <= 1'b0;
			12'd2496: q <= 1'b0;
			12'd2497: q <= 1'b0;
			12'd2498: q <= 1'b0;
			12'd2499: q <= 1'b0;
			12'd2500: q <= 1'b0;
			12'd2501: q <= 1'b0;
			12'd2502: q <= 1'b0;
			12'd2503: q <= 1'b0;
			12'd2504: q <= 1'b0;
			12'd2505: q <= 1'b0;
			12'd2506: q <= 1'b0;
			12'd2507: q <= 1'b0;
			12'd2508: q <= 1'b0;
			12'd2509: q <= 1'b0;
			12'd2510: q <= 1'b0;
			12'd2511: q <= 1'b0;
			12'd2512: q <= 1'b0;
			12'd2513: q <= 1'b0;
			12'd2514: q <= 1'b0;
			12'd2515: q <= 1'b0;
			12'd2516: q <= 1'b0;
			12'd2517: q <= 1'b0;
			12'd2518: q <= 1'b0;
			12'd2519: q <= 1'b0;
			12'd2520: q <= 1'b0;
			12'd2521: q <= 1'b0;
			12'd2522: q <= 1'b0;
			12'd2523: q <= 1'b0;
			12'd2524: q <= 1'b0;
			12'd2525: q <= 1'b0;
			12'd2526: q <= 1'b0;
			12'd2527: q <= 1'b0;
			12'd2528: q <= 1'b0;
			12'd2529: q <= 1'b0;
			12'd2530: q <= 1'b0;
			12'd2531: q <= 1'b0;
			12'd2532: q <= 1'b0;
			12'd2533: q <= 1'b0;
			12'd2534: q <= 1'b0;
			12'd2535: q <= 1'b0;
			12'd2536: q <= 1'b0;
			12'd2537: q <= 1'b0;
			12'd2538: q <= 1'b0;
			12'd2539: q <= 1'b0;
			12'd2540: q <= 1'b0;
			12'd2541: q <= 1'b0;
			12'd2542: q <= 1'b0;
			12'd2543: q <= 1'b0;
			12'd2544: q <= 1'b0;
			12'd2545: q <= 1'b0;
			12'd2546: q <= 1'b0;
			12'd2547: q <= 1'b0;
			12'd2548: q <= 1'b0;
			12'd2549: q <= 1'b0;
			12'd2550: q <= 1'b0;
			12'd2551: q <= 1'b0;
			12'd2552: q <= 1'b0;
			12'd2553: q <= 1'b0;
			12'd2554: q <= 1'b0;
			12'd2555: q <= 1'b0;
			12'd2556: q <= 1'b0;
			12'd2557: q <= 1'b0;
			12'd2558: q <= 1'b0;
			12'd2559: q <= 1'b0;
			12'd2560: q <= 1'b0;
			12'd2561: q <= 1'b0;
			12'd2562: q <= 1'b0;
			12'd2563: q <= 1'b0;
			12'd2564: q <= 1'b0;
			12'd2565: q <= 1'b0;
			12'd2566: q <= 1'b0;
			12'd2567: q <= 1'b0;
			12'd2568: q <= 1'b0;
			12'd2569: q <= 1'b0;
			12'd2570: q <= 1'b0;
			12'd2571: q <= 1'b0;
			12'd2572: q <= 1'b0;
			12'd2573: q <= 1'b0;
			12'd2574: q <= 1'b0;
			12'd2575: q <= 1'b0;
			12'd2576: q <= 1'b0;
			12'd2577: q <= 1'b0;
			12'd2578: q <= 1'b0;
			12'd2579: q <= 1'b0;
			12'd2580: q <= 1'b0;
			12'd2581: q <= 1'b0;
			12'd2582: q <= 1'b0;
			12'd2583: q <= 1'b0;
			12'd2584: q <= 1'b0;
			12'd2585: q <= 1'b0;
			12'd2586: q <= 1'b0;
			12'd2587: q <= 1'b0;
			12'd2588: q <= 1'b0;
			12'd2589: q <= 1'b0;
			12'd2590: q <= 1'b0;
			12'd2591: q <= 1'b0;
			12'd2592: q <= 1'b0;
			12'd2593: q <= 1'b0;
			12'd2594: q <= 1'b0;
			12'd2595: q <= 1'b0;
			12'd2596: q <= 1'b0;
			12'd2597: q <= 1'b0;
			12'd2598: q <= 1'b0;
			12'd2599: q <= 1'b0;
			12'd2600: q <= 1'b0;
			12'd2601: q <= 1'b0;
			12'd2602: q <= 1'b0;
			12'd2603: q <= 1'b0;
			12'd2604: q <= 1'b0;
			12'd2605: q <= 1'b0;
			12'd2606: q <= 1'b0;
			12'd2607: q <= 1'b0;
			12'd2608: q <= 1'b0;
			12'd2609: q <= 1'b0;
			12'd2610: q <= 1'b0;
			12'd2611: q <= 1'b0;
			12'd2612: q <= 1'b0;
			12'd2613: q <= 1'b0;
			12'd2614: q <= 1'b0;
			12'd2615: q <= 1'b0;
			12'd2616: q <= 1'b0;
			12'd2617: q <= 1'b0;
			12'd2618: q <= 1'b0;
			12'd2619: q <= 1'b0;
			12'd2620: q <= 1'b0;
			12'd2621: q <= 1'b0;
			12'd2622: q <= 1'b0;
			12'd2623: q <= 1'b0;
			12'd2624: q <= 1'b0;
			12'd2625: q <= 1'b0;
			12'd2626: q <= 1'b0;
			12'd2627: q <= 1'b0;
			12'd2628: q <= 1'b0;
			12'd2629: q <= 1'b0;
			12'd2630: q <= 1'b0;
			12'd2631: q <= 1'b0;
			12'd2632: q <= 1'b0;
			12'd2633: q <= 1'b0;
			12'd2634: q <= 1'b0;
			12'd2635: q <= 1'b0;
			12'd2636: q <= 1'b0;
			12'd2637: q <= 1'b0;
			12'd2638: q <= 1'b0;
			12'd2639: q <= 1'b0;
			12'd2640: q <= 1'b0;
			12'd2641: q <= 1'b0;
			12'd2642: q <= 1'b0;
			12'd2643: q <= 1'b0;
			12'd2644: q <= 1'b0;
			12'd2645: q <= 1'b0;
			12'd2646: q <= 1'b0;
			12'd2647: q <= 1'b0;
			12'd2648: q <= 1'b0;
			12'd2649: q <= 1'b0;
			12'd2650: q <= 1'b0;
			12'd2651: q <= 1'b0;
			12'd2652: q <= 1'b0;
			12'd2653: q <= 1'b0;
			12'd2654: q <= 1'b0;
			12'd2655: q <= 1'b0;
			12'd2656: q <= 1'b0;
			12'd2657: q <= 1'b0;
			12'd2658: q <= 1'b0;
			12'd2659: q <= 1'b0;
			12'd2660: q <= 1'b0;
			12'd2661: q <= 1'b0;
			12'd2662: q <= 1'b0;
			12'd2663: q <= 1'b0;
			12'd2664: q <= 1'b0;
			12'd2665: q <= 1'b0;
			12'd2666: q <= 1'b0;
			12'd2667: q <= 1'b0;
			12'd2668: q <= 1'b0;
			12'd2669: q <= 1'b0;
			12'd2670: q <= 1'b0;
			12'd2671: q <= 1'b0;
			12'd2672: q <= 1'b0;
			12'd2673: q <= 1'b0;
			12'd2674: q <= 1'b0;
			12'd2675: q <= 1'b0;
			12'd2676: q <= 1'b0;
			12'd2677: q <= 1'b0;
			12'd2678: q <= 1'b0;
			12'd2679: q <= 1'b0;
			12'd2680: q <= 1'b0;
			12'd2681: q <= 1'b0;
			12'd2682: q <= 1'b0;
			12'd2683: q <= 1'b0;
			12'd2684: q <= 1'b0;
			12'd2685: q <= 1'b0;
			12'd2686: q <= 1'b0;
			12'd2687: q <= 1'b0;
			12'd2688: q <= 1'b0;
			12'd2689: q <= 1'b0;
			12'd2690: q <= 1'b0;
			12'd2691: q <= 1'b0;
			12'd2692: q <= 1'b0;
			12'd2693: q <= 1'b0;
			12'd2694: q <= 1'b0;
			12'd2695: q <= 1'b0;
			12'd2696: q <= 1'b0;
			12'd2697: q <= 1'b0;
			12'd2698: q <= 1'b0;
			12'd2699: q <= 1'b0;
			12'd2700: q <= 1'b0;
			12'd2701: q <= 1'b0;
			12'd2702: q <= 1'b0;
			12'd2703: q <= 1'b0;
			12'd2704: q <= 1'b0;
			12'd2705: q <= 1'b0;
			12'd2706: q <= 1'b0;
			12'd2707: q <= 1'b0;
			12'd2708: q <= 1'b0;
			12'd2709: q <= 1'b0;
			12'd2710: q <= 1'b0;
			12'd2711: q <= 1'b0;
			12'd2712: q <= 1'b0;
			12'd2713: q <= 1'b0;
			12'd2714: q <= 1'b0;
			12'd2715: q <= 1'b0;
			12'd2716: q <= 1'b0;
			12'd2717: q <= 1'b0;
			12'd2718: q <= 1'b0;
			12'd2719: q <= 1'b0;
			12'd2720: q <= 1'b0;
			12'd2721: q <= 1'b0;
			12'd2722: q <= 1'b0;
			12'd2723: q <= 1'b0;
			12'd2724: q <= 1'b0;
			12'd2725: q <= 1'b0;
			12'd2726: q <= 1'b0;
			12'd2727: q <= 1'b0;
			12'd2728: q <= 1'b0;
			12'd2729: q <= 1'b0;
			12'd2730: q <= 1'b0;
			12'd2731: q <= 1'b0;
			12'd2732: q <= 1'b0;
			12'd2733: q <= 1'b0;
			12'd2734: q <= 1'b0;
			12'd2735: q <= 1'b0;
			12'd2736: q <= 1'b0;
			12'd2737: q <= 1'b0;
			12'd2738: q <= 1'b0;
			12'd2739: q <= 1'b0;
			12'd2740: q <= 1'b0;
			12'd2741: q <= 1'b0;
			12'd2742: q <= 1'b0;
			12'd2743: q <= 1'b0;
			12'd2744: q <= 1'b0;
			12'd2745: q <= 1'b0;
			12'd2746: q <= 1'b0;
			12'd2747: q <= 1'b0;
			12'd2748: q <= 1'b0;
			12'd2749: q <= 1'b0;
			12'd2750: q <= 1'b0;
			12'd2751: q <= 1'b0;
			12'd2752: q <= 1'b0;
			12'd2753: q <= 1'b0;
			12'd2754: q <= 1'b0;
			12'd2755: q <= 1'b0;
			12'd2756: q <= 1'b0;
			12'd2757: q <= 1'b0;
			12'd2758: q <= 1'b0;
			12'd2759: q <= 1'b0;
			12'd2760: q <= 1'b0;
			12'd2761: q <= 1'b0;
			12'd2762: q <= 1'b0;
			12'd2763: q <= 1'b0;
			12'd2764: q <= 1'b0;
			12'd2765: q <= 1'b0;
			12'd2766: q <= 1'b0;
			12'd2767: q <= 1'b0;
			12'd2768: q <= 1'b0;
			12'd2769: q <= 1'b0;
			12'd2770: q <= 1'b0;
			12'd2771: q <= 1'b0;
			12'd2772: q <= 1'b0;
			12'd2773: q <= 1'b0;
			12'd2774: q <= 1'b0;
			12'd2775: q <= 1'b0;
			12'd2776: q <= 1'b0;
			12'd2777: q <= 1'b0;
			12'd2778: q <= 1'b0;
			12'd2779: q <= 1'b0;
			12'd2780: q <= 1'b0;
			12'd2781: q <= 1'b0;
			12'd2782: q <= 1'b0;
			12'd2783: q <= 1'b0;
			12'd2784: q <= 1'b0;
			12'd2785: q <= 1'b0;
			12'd2786: q <= 1'b0;
			12'd2787: q <= 1'b0;
			12'd2788: q <= 1'b0;
			12'd2789: q <= 1'b0;
			12'd2790: q <= 1'b0;
			12'd2791: q <= 1'b0;
			12'd2792: q <= 1'b0;
			12'd2793: q <= 1'b0;
			12'd2794: q <= 1'b0;
			12'd2795: q <= 1'b0;
			12'd2796: q <= 1'b0;
			12'd2797: q <= 1'b0;
			12'd2798: q <= 1'b0;
			12'd2799: q <= 1'b0;
			12'd2800: q <= 1'b0;
			12'd2801: q <= 1'b0;
			12'd2802: q <= 1'b0;
			12'd2803: q <= 1'b0;
			12'd2804: q <= 1'b0;
			12'd2805: q <= 1'b0;
			12'd2806: q <= 1'b0;
			12'd2807: q <= 1'b0;
			12'd2808: q <= 1'b0;
			12'd2809: q <= 1'b0;
			12'd2810: q <= 1'b0;
			12'd2811: q <= 1'b0;
			12'd2812: q <= 1'b0;
			12'd2813: q <= 1'b0;
			12'd2814: q <= 1'b0;
			12'd2815: q <= 1'b0;
			12'd2816: q <= 1'b0;
			12'd2817: q <= 1'b0;
			12'd2818: q <= 1'b0;
			12'd2819: q <= 1'b0;
			12'd2820: q <= 1'b0;
			12'd2821: q <= 1'b0;
			12'd2822: q <= 1'b0;
			12'd2823: q <= 1'b0;
			12'd2824: q <= 1'b0;
			12'd2825: q <= 1'b0;
			12'd2826: q <= 1'b0;
			12'd2827: q <= 1'b0;
			12'd2828: q <= 1'b0;
			12'd2829: q <= 1'b0;
			12'd2830: q <= 1'b0;
			12'd2831: q <= 1'b0;
			12'd2832: q <= 1'b0;
			12'd2833: q <= 1'b0;
			12'd2834: q <= 1'b0;
			12'd2835: q <= 1'b1;
			12'd2836: q <= 1'b1;
			12'd2837: q <= 1'b1;
			12'd2838: q <= 1'b1;
			12'd2839: q <= 1'b1;
			12'd2840: q <= 1'b1;
			12'd2841: q <= 1'b1;
			12'd2842: q <= 1'b1;
			12'd2843: q <= 1'b1;
			12'd2844: q <= 1'b1;
			12'd2845: q <= 1'b1;
			12'd2846: q <= 1'b1;
			12'd2847: q <= 1'b1;
			12'd2848: q <= 1'b1;
			12'd2849: q <= 1'b1;
			12'd2850: q <= 1'b0;
			12'd2851: q <= 1'b0;
			12'd2852: q <= 1'b0;
			12'd2853: q <= 1'b0;
			12'd2854: q <= 1'b0;
			12'd2855: q <= 1'b0;
			12'd2856: q <= 1'b0;
			12'd2857: q <= 1'b0;
			12'd2858: q <= 1'b0;
			12'd2859: q <= 1'b0;
			12'd2860: q <= 1'b0;
			12'd2861: q <= 1'b0;
			12'd2862: q <= 1'b0;
			12'd2863: q <= 1'b0;
			12'd2864: q <= 1'b0;
			12'd2865: q <= 1'b1;
			12'd2866: q <= 1'b1;
			12'd2867: q <= 1'b1;
			12'd2868: q <= 1'b1;
			12'd2869: q <= 1'b1;
			12'd2870: q <= 1'b1;
			12'd2871: q <= 1'b1;
			12'd2872: q <= 1'b1;
			12'd2873: q <= 1'b1;
			12'd2874: q <= 1'b1;
			12'd2875: q <= 1'b1;
			12'd2876: q <= 1'b1;
			12'd2877: q <= 1'b1;
			12'd2878: q <= 1'b1;
			12'd2879: q <= 1'b1;
			12'd2880: q <= 1'b1;
			12'd2881: q <= 1'b1;
			12'd2882: q <= 1'b1;
			12'd2883: q <= 1'b1;
			12'd2884: q <= 1'b1;
			12'd2885: q <= 1'b1;
			12'd2886: q <= 1'b1;
			12'd2887: q <= 1'b1;
			12'd2888: q <= 1'b1;
			12'd2889: q <= 1'b1;
			12'd2890: q <= 1'b0;
			12'd2891: q <= 1'b0;
			12'd2892: q <= 1'b0;
			12'd2893: q <= 1'b0;
			12'd2894: q <= 1'b0;
			12'd2895: q <= 1'b0;
			12'd2896: q <= 1'b0;
			12'd2897: q <= 1'b0;
			12'd2898: q <= 1'b0;
			12'd2899: q <= 1'b0;
			12'd2900: q <= 1'b0;
			12'd2901: q <= 1'b0;
			12'd2902: q <= 1'b0;
			12'd2903: q <= 1'b0;
			12'd2904: q <= 1'b0;
			12'd2905: q <= 1'b1;
			12'd2906: q <= 1'b1;
			12'd2907: q <= 1'b1;
			12'd2908: q <= 1'b1;
			12'd2909: q <= 1'b1;
			12'd2910: q <= 1'b1;
			12'd2911: q <= 1'b1;
			12'd2912: q <= 1'b1;
			12'd2913: q <= 1'b1;
			12'd2914: q <= 1'b1;
			12'd2915: q <= 1'b1;
			12'd2916: q <= 1'b1;
			12'd2917: q <= 1'b1;
			12'd2918: q <= 1'b1;
			12'd2919: q <= 1'b1;
			12'd2920: q <= 1'b1;
			12'd2921: q <= 1'b1;
			12'd2922: q <= 1'b1;
			12'd2923: q <= 1'b1;
			12'd2924: q <= 1'b1;
			12'd2925: q <= 1'b1;
			12'd2926: q <= 1'b1;
			12'd2927: q <= 1'b1;
			12'd2928: q <= 1'b1;
			12'd2929: q <= 1'b1;
			12'd2930: q <= 1'b0;
			12'd2931: q <= 1'b0;
			12'd2932: q <= 1'b0;
			12'd2933: q <= 1'b0;
			12'd2934: q <= 1'b0;
			12'd2935: q <= 1'b0;
			12'd2936: q <= 1'b0;
			12'd2937: q <= 1'b0;
			12'd2938: q <= 1'b0;
			12'd2939: q <= 1'b0;
			12'd2940: q <= 1'b0;
			12'd2941: q <= 1'b0;
			12'd2942: q <= 1'b0;
			12'd2943: q <= 1'b0;
			12'd2944: q <= 1'b0;
			12'd2945: q <= 1'b0;
			12'd2946: q <= 1'b1;
			12'd2947: q <= 1'b1;
			12'd2948: q <= 1'b1;
			12'd2949: q <= 1'b1;
			12'd2950: q <= 1'b1;
			12'd2951: q <= 1'b1;
			12'd2952: q <= 1'b1;
			12'd2953: q <= 1'b1;
			12'd2954: q <= 1'b1;
			12'd2955: q <= 1'b1;
			12'd2956: q <= 1'b1;
			12'd2957: q <= 1'b1;
			12'd2958: q <= 1'b1;
			12'd2959: q <= 1'b1;
			12'd2960: q <= 1'b1;
			12'd2961: q <= 1'b1;
			12'd2962: q <= 1'b1;
			12'd2963: q <= 1'b1;
			12'd2964: q <= 1'b1;
			12'd2965: q <= 1'b1;
			12'd2966: q <= 1'b1;
			12'd2967: q <= 1'b1;
			12'd2968: q <= 1'b1;
			12'd2969: q <= 1'b1;
			12'd2970: q <= 1'b0;
			12'd2971: q <= 1'b0;
			12'd2972: q <= 1'b0;
			12'd2973: q <= 1'b0;
			12'd2974: q <= 1'b0;
			12'd2975: q <= 1'b0;
			12'd2976: q <= 1'b0;
			12'd2977: q <= 1'b0;
			12'd2978: q <= 1'b0;
			12'd2979: q <= 1'b0;
			12'd2980: q <= 1'b0;
			12'd2981: q <= 1'b0;
			12'd2982: q <= 1'b0;
			12'd2983: q <= 1'b0;
			12'd2984: q <= 1'b1;
			12'd2985: q <= 1'b1;
			12'd2986: q <= 1'b1;
			12'd2987: q <= 1'b1;
			12'd2988: q <= 1'b1;
			12'd2989: q <= 1'b1;
			12'd2990: q <= 1'b1;
			12'd2991: q <= 1'b1;
			12'd2992: q <= 1'b1;
			12'd2993: q <= 1'b1;
			12'd2994: q <= 1'b1;
			12'd2995: q <= 1'b1;
			12'd2996: q <= 1'b1;
			12'd2997: q <= 1'b1;
			12'd2998: q <= 1'b1;
			12'd2999: q <= 1'b1;
			12'd3000: q <= 1'b1;
			12'd3001: q <= 1'b1;
			12'd3002: q <= 1'b1;
			12'd3003: q <= 1'b1;
			12'd3004: q <= 1'b1;
			12'd3005: q <= 1'b1;
			12'd3006: q <= 1'b1;
			12'd3007: q <= 1'b1;
			12'd3008: q <= 1'b1;
			12'd3009: q <= 1'b1;
			12'd3010: q <= 1'b0;
			12'd3011: q <= 1'b0;
			12'd3012: q <= 1'b0;
			12'd3013: q <= 1'b0;
			12'd3014: q <= 1'b0;
			12'd3015: q <= 1'b0;
			12'd3016: q <= 1'b0;
			12'd3017: q <= 1'b0;
			12'd3018: q <= 1'b0;
			12'd3019: q <= 1'b0;
			12'd3020: q <= 1'b0;
			12'd3021: q <= 1'b0;
			12'd3022: q <= 1'b0;
			12'd3023: q <= 1'b0;
			12'd3024: q <= 1'b1;
			12'd3025: q <= 1'b1;
			12'd3026: q <= 1'b1;
			12'd3027: q <= 1'b1;
			12'd3028: q <= 1'b1;
			12'd3029: q <= 1'b1;
			12'd3030: q <= 1'b1;
			12'd3031: q <= 1'b1;
			12'd3032: q <= 1'b1;
			12'd3033: q <= 1'b1;
			12'd3034: q <= 1'b1;
			12'd3035: q <= 1'b1;
			12'd3036: q <= 1'b1;
			12'd3037: q <= 1'b1;
			12'd3038: q <= 1'b1;
			12'd3039: q <= 1'b1;
			12'd3040: q <= 1'b1;
			12'd3041: q <= 1'b1;
			12'd3042: q <= 1'b1;
			12'd3043: q <= 1'b1;
			12'd3044: q <= 1'b1;
			12'd3045: q <= 1'b1;
			12'd3046: q <= 1'b1;
			12'd3047: q <= 1'b1;
			12'd3048: q <= 1'b1;
			12'd3049: q <= 1'b1;
			12'd3050: q <= 1'b0;
			12'd3051: q <= 1'b0;
			12'd3052: q <= 1'b0;
			12'd3053: q <= 1'b0;
			12'd3054: q <= 1'b0;
			12'd3055: q <= 1'b0;
			12'd3056: q <= 1'b0;
			12'd3057: q <= 1'b0;
			12'd3058: q <= 1'b0;
			12'd3059: q <= 1'b0;
			12'd3060: q <= 1'b0;
			12'd3061: q <= 1'b0;
			12'd3062: q <= 1'b0;
			12'd3063: q <= 1'b1;
			12'd3064: q <= 1'b1;
			12'd3065: q <= 1'b1;
			12'd3066: q <= 1'b1;
			12'd3067: q <= 1'b1;
			12'd3068: q <= 1'b1;
			12'd3069: q <= 1'b1;
			12'd3070: q <= 1'b1;
			12'd3071: q <= 1'b1;
			12'd3072: q <= 1'b1;
			12'd3073: q <= 1'b1;
			12'd3074: q <= 1'b1;
			12'd3075: q <= 1'b1;
			12'd3076: q <= 1'b1;
			12'd3077: q <= 1'b1;
			12'd3078: q <= 1'b1;
			12'd3079: q <= 1'b1;
			12'd3080: q <= 1'b1;
			12'd3081: q <= 1'b1;
			12'd3082: q <= 1'b1;
			12'd3083: q <= 1'b1;
			12'd3084: q <= 1'b1;
			12'd3085: q <= 1'b1;
			12'd3086: q <= 1'b1;
			12'd3087: q <= 1'b1;
			12'd3088: q <= 1'b1;
			12'd3089: q <= 1'b1;
			12'd3090: q <= 1'b0;
			12'd3091: q <= 1'b0;
			12'd3092: q <= 1'b0;
			12'd3093: q <= 1'b0;
			12'd3094: q <= 1'b0;
			12'd3095: q <= 1'b0;
			12'd3096: q <= 1'b0;
			12'd3097: q <= 1'b0;
			12'd3098: q <= 1'b0;
			12'd3099: q <= 1'b0;
			12'd3100: q <= 1'b0;
			12'd3101: q <= 1'b0;
			12'd3102: q <= 1'b0;
			12'd3103: q <= 1'b1;
			12'd3104: q <= 1'b1;
			12'd3105: q <= 1'b1;
			12'd3106: q <= 1'b1;
			12'd3107: q <= 1'b1;
			12'd3108: q <= 1'b1;
			12'd3109: q <= 1'b1;
			12'd3110: q <= 1'b1;
			12'd3111: q <= 1'b1;
			12'd3112: q <= 1'b1;
			12'd3113: q <= 1'b1;
			12'd3114: q <= 1'b1;
			12'd3115: q <= 1'b1;
			12'd3116: q <= 1'b1;
			12'd3117: q <= 1'b1;
			12'd3118: q <= 1'b1;
			12'd3119: q <= 1'b1;
			12'd3120: q <= 1'b1;
			12'd3121: q <= 1'b1;
			12'd3122: q <= 1'b1;
			12'd3123: q <= 1'b1;
			12'd3124: q <= 1'b1;
			12'd3125: q <= 1'b1;
			12'd3126: q <= 1'b1;
			12'd3127: q <= 1'b1;
			12'd3128: q <= 1'b1;
			12'd3129: q <= 1'b1;
			12'd3130: q <= 1'b0;
			12'd3131: q <= 1'b0;
			12'd3132: q <= 1'b0;
			12'd3133: q <= 1'b0;
			12'd3134: q <= 1'b0;
			12'd3135: q <= 1'b0;
			12'd3136: q <= 1'b0;
			12'd3137: q <= 1'b0;
			12'd3138: q <= 1'b0;
			12'd3139: q <= 1'b0;
			12'd3140: q <= 1'b0;
			12'd3141: q <= 1'b0;
			12'd3142: q <= 1'b0;
			12'd3143: q <= 1'b1;
			12'd3144: q <= 1'b1;
			12'd3145: q <= 1'b1;
			12'd3146: q <= 1'b1;
			12'd3147: q <= 1'b1;
			12'd3148: q <= 1'b1;
			12'd3149: q <= 1'b1;
			12'd3150: q <= 1'b1;
			12'd3151: q <= 1'b1;
			12'd3152: q <= 1'b1;
			12'd3153: q <= 1'b1;
			12'd3154: q <= 1'b1;
			12'd3155: q <= 1'b1;
			12'd3156: q <= 1'b1;
			12'd3157: q <= 1'b1;
			12'd3158: q <= 1'b1;
			12'd3159: q <= 1'b1;
			12'd3160: q <= 1'b1;
			12'd3161: q <= 1'b1;
			12'd3162: q <= 1'b1;
			12'd3163: q <= 1'b1;
			12'd3164: q <= 1'b1;
			12'd3165: q <= 1'b1;
			12'd3166: q <= 1'b1;
			12'd3167: q <= 1'b1;
			12'd3168: q <= 1'b1;
			12'd3169: q <= 1'b1;
			12'd3170: q <= 1'b1;
			12'd3171: q <= 1'b0;
			12'd3172: q <= 1'b0;
			12'd3173: q <= 1'b0;
			12'd3174: q <= 1'b0;
			12'd3175: q <= 1'b0;
			12'd3176: q <= 1'b0;
			12'd3177: q <= 1'b0;
			12'd3178: q <= 1'b0;
			12'd3179: q <= 1'b0;
			12'd3180: q <= 1'b0;
			12'd3181: q <= 1'b0;
			12'd3182: q <= 1'b0;
			12'd3183: q <= 1'b1;
			12'd3184: q <= 1'b1;
			12'd3185: q <= 1'b1;
			12'd3186: q <= 1'b1;
			12'd3187: q <= 1'b1;
			12'd3188: q <= 1'b1;
			12'd3189: q <= 1'b1;
			12'd3190: q <= 1'b1;
			12'd3191: q <= 1'b1;
			12'd3192: q <= 1'b1;
			12'd3193: q <= 1'b1;
			12'd3194: q <= 1'b1;
			12'd3195: q <= 1'b1;
			12'd3196: q <= 1'b1;
			12'd3197: q <= 1'b1;
			12'd3198: q <= 1'b1;
			12'd3199: q <= 1'b1;
			12'd3200: q <= 1'b1;
			12'd3201: q <= 1'b1;
			12'd3202: q <= 1'b1;
			12'd3203: q <= 1'b1;
			12'd3204: q <= 1'b1;
			12'd3205: q <= 1'b1;
			12'd3206: q <= 1'b1;
			12'd3207: q <= 1'b1;
			12'd3208: q <= 1'b1;
			12'd3209: q <= 1'b1;
			12'd3210: q <= 1'b1;
			12'd3211: q <= 1'b1;
			12'd3212: q <= 1'b0;
			12'd3213: q <= 1'b0;
			12'd3214: q <= 1'b0;
			12'd3215: q <= 1'b0;
			12'd3216: q <= 1'b0;
			12'd3217: q <= 1'b0;
			12'd3218: q <= 1'b0;
			12'd3219: q <= 1'b0;
			12'd3220: q <= 1'b0;
			12'd3221: q <= 1'b0;
			12'd3222: q <= 1'b0;
			12'd3223: q <= 1'b1;
			12'd3224: q <= 1'b1;
			12'd3225: q <= 1'b1;
			12'd3226: q <= 1'b1;
			12'd3227: q <= 1'b1;
			12'd3228: q <= 1'b1;
			12'd3229: q <= 1'b1;
			12'd3230: q <= 1'b1;
			12'd3231: q <= 1'b1;
			12'd3232: q <= 1'b1;
			12'd3233: q <= 1'b1;
			12'd3234: q <= 1'b1;
			12'd3235: q <= 1'b1;
			12'd3236: q <= 1'b1;
			12'd3237: q <= 1'b1;
			12'd3238: q <= 1'b1;
			12'd3239: q <= 1'b1;
			12'd3240: q <= 1'b1;
			12'd3241: q <= 1'b1;
			12'd3242: q <= 1'b1;
			12'd3243: q <= 1'b1;
			12'd3244: q <= 1'b1;
			12'd3245: q <= 1'b1;
			12'd3246: q <= 1'b1;
			12'd3247: q <= 1'b1;
			12'd3248: q <= 1'b1;
			12'd3249: q <= 1'b1;
			12'd3250: q <= 1'b1;
			12'd3251: q <= 1'b1;
			12'd3252: q <= 1'b1;
			12'd3253: q <= 1'b1;
			12'd3254: q <= 1'b0;
			12'd3255: q <= 1'b0;
			12'd3256: q <= 1'b0;
			12'd3257: q <= 1'b0;
			12'd3258: q <= 1'b0;
			12'd3259: q <= 1'b0;
			12'd3260: q <= 1'b0;
			12'd3261: q <= 1'b0;
			12'd3262: q <= 1'b0;
			12'd3263: q <= 1'b1;
			12'd3264: q <= 1'b1;
			12'd3265: q <= 1'b1;
			12'd3266: q <= 1'b1;
			12'd3267: q <= 1'b1;
			12'd3268: q <= 1'b1;
			12'd3269: q <= 1'b1;
			12'd3270: q <= 1'b1;
			12'd3271: q <= 1'b1;
			12'd3272: q <= 1'b1;
			12'd3273: q <= 1'b1;
			12'd3274: q <= 1'b1;
			12'd3275: q <= 1'b1;
			12'd3276: q <= 1'b1;
			12'd3277: q <= 1'b1;
			12'd3278: q <= 1'b1;
			12'd3279: q <= 1'b1;
			12'd3280: q <= 1'b1;
			12'd3281: q <= 1'b1;
			12'd3282: q <= 1'b1;
			12'd3283: q <= 1'b1;
			12'd3284: q <= 1'b1;
			12'd3285: q <= 1'b1;
			12'd3286: q <= 1'b1;
			12'd3287: q <= 1'b1;
			12'd3288: q <= 1'b1;
			12'd3289: q <= 1'b1;
			12'd3290: q <= 1'b1;
			12'd3291: q <= 1'b1;
			12'd3292: q <= 1'b1;
			12'd3293: q <= 1'b1;
			12'd3294: q <= 1'b1;
			12'd3295: q <= 1'b0;
			12'd3296: q <= 1'b0;
			12'd3297: q <= 1'b0;
			12'd3298: q <= 1'b0;
			12'd3299: q <= 1'b0;
			12'd3300: q <= 1'b0;
			12'd3301: q <= 1'b0;
			12'd3302: q <= 1'b0;
			12'd3303: q <= 1'b1;
			12'd3304: q <= 1'b1;
			12'd3305: q <= 1'b1;
			12'd3306: q <= 1'b1;
			12'd3307: q <= 1'b1;
			12'd3308: q <= 1'b1;
			12'd3309: q <= 1'b1;
			12'd3310: q <= 1'b1;
			12'd3311: q <= 1'b1;
			12'd3312: q <= 1'b1;
			12'd3313: q <= 1'b1;
			12'd3314: q <= 1'b1;
			12'd3315: q <= 1'b1;
			12'd3316: q <= 1'b1;
			12'd3317: q <= 1'b1;
			12'd3318: q <= 1'b1;
			12'd3319: q <= 1'b1;
			12'd3320: q <= 1'b1;
			12'd3321: q <= 1'b1;
			12'd3322: q <= 1'b1;
			12'd3323: q <= 1'b1;
			12'd3324: q <= 1'b1;
			12'd3325: q <= 1'b1;
			12'd3326: q <= 1'b1;
			12'd3327: q <= 1'b1;
			12'd3328: q <= 1'b1;
			12'd3329: q <= 1'b1;
			12'd3330: q <= 1'b1;
			12'd3331: q <= 1'b1;
			12'd3332: q <= 1'b1;
			12'd3333: q <= 1'b1;
			12'd3334: q <= 1'b1;
			12'd3335: q <= 1'b1;
			12'd3336: q <= 1'b0;
			12'd3337: q <= 1'b0;
			12'd3338: q <= 1'b0;
			12'd3339: q <= 1'b0;
			12'd3340: q <= 1'b0;
			12'd3341: q <= 1'b0;
			12'd3342: q <= 1'b0;
			12'd3343: q <= 1'b1;
			12'd3344: q <= 1'b1;
			12'd3345: q <= 1'b1;
			12'd3346: q <= 1'b1;
			12'd3347: q <= 1'b1;
			12'd3348: q <= 1'b1;
			12'd3349: q <= 1'b1;
			12'd3350: q <= 1'b1;
			12'd3351: q <= 1'b1;
			12'd3352: q <= 1'b1;
			12'd3353: q <= 1'b1;
			12'd3354: q <= 1'b1;
			12'd3355: q <= 1'b1;
			12'd3356: q <= 1'b1;
			12'd3357: q <= 1'b1;
			12'd3358: q <= 1'b1;
			12'd3359: q <= 1'b1;
			12'd3360: q <= 1'b1;
			12'd3361: q <= 1'b1;
			12'd3362: q <= 1'b1;
			12'd3363: q <= 1'b1;
			12'd3364: q <= 1'b1;
			12'd3365: q <= 1'b1;
			12'd3366: q <= 1'b1;
			12'd3367: q <= 1'b1;
			12'd3368: q <= 1'b1;
			12'd3369: q <= 1'b1;
			12'd3370: q <= 1'b1;
			12'd3371: q <= 1'b1;
			12'd3372: q <= 1'b1;
			12'd3373: q <= 1'b1;
			12'd3374: q <= 1'b1;
			12'd3375: q <= 1'b1;
			12'd3376: q <= 1'b0;
			12'd3377: q <= 1'b0;
			12'd3378: q <= 1'b0;
			12'd3379: q <= 1'b0;
			12'd3380: q <= 1'b0;
			12'd3381: q <= 1'b0;
			12'd3382: q <= 1'b1;
			12'd3383: q <= 1'b1;
			12'd3384: q <= 1'b1;
			12'd3385: q <= 1'b1;
			12'd3386: q <= 1'b1;
			12'd3387: q <= 1'b1;
			12'd3388: q <= 1'b1;
			12'd3389: q <= 1'b1;
			12'd3390: q <= 1'b1;
			12'd3391: q <= 1'b1;
			12'd3392: q <= 1'b1;
			12'd3393: q <= 1'b1;
			12'd3394: q <= 1'b1;
			12'd3395: q <= 1'b1;
			12'd3396: q <= 1'b1;
			12'd3397: q <= 1'b1;
			12'd3398: q <= 1'b1;
			12'd3399: q <= 1'b1;
			12'd3400: q <= 1'b1;
			12'd3401: q <= 1'b1;
			12'd3402: q <= 1'b1;
			12'd3403: q <= 1'b1;
			12'd3404: q <= 1'b1;
			12'd3405: q <= 1'b1;
			12'd3406: q <= 1'b1;
			12'd3407: q <= 1'b1;
			12'd3408: q <= 1'b1;
			12'd3409: q <= 1'b1;
			12'd3410: q <= 1'b1;
			12'd3411: q <= 1'b1;
			12'd3412: q <= 1'b1;
			12'd3413: q <= 1'b1;
			12'd3414: q <= 1'b1;
			12'd3415: q <= 1'b1;
			12'd3416: q <= 1'b1;
			12'd3417: q <= 1'b0;
			12'd3418: q <= 1'b0;
			12'd3419: q <= 1'b0;
			12'd3420: q <= 1'b0;
			12'd3421: q <= 1'b0;
			12'd3422: q <= 1'b1;
			12'd3423: q <= 1'b1;
			12'd3424: q <= 1'b1;
			12'd3425: q <= 1'b1;
			12'd3426: q <= 1'b1;
			12'd3427: q <= 1'b1;
			12'd3428: q <= 1'b1;
			12'd3429: q <= 1'b1;
			12'd3430: q <= 1'b1;
			12'd3431: q <= 1'b1;
			12'd3432: q <= 1'b1;
			12'd3433: q <= 1'b1;
			12'd3434: q <= 1'b1;
			12'd3435: q <= 1'b1;
			12'd3436: q <= 1'b1;
			12'd3437: q <= 1'b1;
			12'd3438: q <= 1'b1;
			12'd3439: q <= 1'b1;
			12'd3440: q <= 1'b1;
			12'd3441: q <= 1'b1;
			12'd3442: q <= 1'b1;
			12'd3443: q <= 1'b1;
			12'd3444: q <= 1'b1;
			12'd3445: q <= 1'b1;
			12'd3446: q <= 1'b1;
			12'd3447: q <= 1'b1;
			12'd3448: q <= 1'b1;
			12'd3449: q <= 1'b1;
			12'd3450: q <= 1'b1;
			12'd3451: q <= 1'b1;
			12'd3452: q <= 1'b1;
			12'd3453: q <= 1'b1;
			12'd3454: q <= 1'b1;
			12'd3455: q <= 1'b1;
			12'd3456: q <= 1'b0;
			12'd3457: q <= 1'b0;
			12'd3458: q <= 1'b0;
			12'd3459: q <= 1'b0;
			12'd3460: q <= 1'b0;
			12'd3461: q <= 1'b0;
			12'd3462: q <= 1'b0;
			12'd3463: q <= 1'b1;
			12'd3464: q <= 1'b1;
			12'd3465: q <= 1'b1;
			12'd3466: q <= 1'b1;
			12'd3467: q <= 1'b1;
			12'd3468: q <= 1'b1;
			12'd3469: q <= 1'b1;
			12'd3470: q <= 1'b1;
			12'd3471: q <= 1'b1;
			12'd3472: q <= 1'b1;
			12'd3473: q <= 1'b1;
			12'd3474: q <= 1'b1;
			12'd3475: q <= 1'b1;
			12'd3476: q <= 1'b1;
			12'd3477: q <= 1'b1;
			12'd3478: q <= 1'b1;
			12'd3479: q <= 1'b1;
			12'd3480: q <= 1'b1;
			12'd3481: q <= 1'b1;
			12'd3482: q <= 1'b1;
			12'd3483: q <= 1'b1;
			12'd3484: q <= 1'b1;
			12'd3485: q <= 1'b1;
			12'd3486: q <= 1'b1;
			12'd3487: q <= 1'b1;
			12'd3488: q <= 1'b1;
			12'd3489: q <= 1'b1;
			12'd3490: q <= 1'b1;
			12'd3491: q <= 1'b1;
			12'd3492: q <= 1'b1;
			12'd3493: q <= 1'b1;
			12'd3494: q <= 1'b1;
			12'd3495: q <= 1'b1;
			12'd3496: q <= 1'b0;
			12'd3497: q <= 1'b0;
			12'd3498: q <= 1'b0;
			12'd3499: q <= 1'b0;
			12'd3500: q <= 1'b0;
			12'd3501: q <= 1'b0;
			12'd3502: q <= 1'b0;
			12'd3503: q <= 1'b1;
			12'd3504: q <= 1'b1;
			12'd3505: q <= 1'b1;
			12'd3506: q <= 1'b1;
			12'd3507: q <= 1'b1;
			12'd3508: q <= 1'b1;
			12'd3509: q <= 1'b1;
			12'd3510: q <= 1'b1;
			12'd3511: q <= 1'b1;
			12'd3512: q <= 1'b1;
			12'd3513: q <= 1'b1;
			12'd3514: q <= 1'b1;
			12'd3515: q <= 1'b1;
			12'd3516: q <= 1'b1;
			12'd3517: q <= 1'b1;
			12'd3518: q <= 1'b1;
			12'd3519: q <= 1'b1;
			12'd3520: q <= 1'b1;
			12'd3521: q <= 1'b1;
			12'd3522: q <= 1'b1;
			12'd3523: q <= 1'b1;
			12'd3524: q <= 1'b1;
			12'd3525: q <= 1'b1;
			12'd3526: q <= 1'b1;
			12'd3527: q <= 1'b1;
			12'd3528: q <= 1'b1;
			12'd3529: q <= 1'b1;
			12'd3530: q <= 1'b1;
			12'd3531: q <= 1'b1;
			12'd3532: q <= 1'b1;
			12'd3533: q <= 1'b1;
			12'd3534: q <= 1'b1;
			12'd3535: q <= 1'b1;
			12'd3536: q <= 1'b1;
			12'd3537: q <= 1'b0;
			12'd3538: q <= 1'b0;
			12'd3539: q <= 1'b0;
			12'd3540: q <= 1'b0;
			12'd3541: q <= 1'b0;
			12'd3542: q <= 1'b0;
			12'd3543: q <= 1'b1;
			12'd3544: q <= 1'b1;
			12'd3545: q <= 1'b1;
			12'd3546: q <= 1'b0;
			12'd3547: q <= 1'b1;
			12'd3548: q <= 1'b1;
			12'd3549: q <= 1'b1;
			12'd3550: q <= 1'b1;
			12'd3551: q <= 1'b1;
			12'd3552: q <= 1'b1;
			12'd3553: q <= 1'b1;
			12'd3554: q <= 1'b1;
			12'd3555: q <= 1'b1;
			12'd3556: q <= 1'b1;
			12'd3557: q <= 1'b1;
			12'd3558: q <= 1'b1;
			12'd3559: q <= 1'b1;
			12'd3560: q <= 1'b1;
			12'd3561: q <= 1'b1;
			12'd3562: q <= 1'b1;
			12'd3563: q <= 1'b1;
			12'd3564: q <= 1'b1;
			12'd3565: q <= 1'b1;
			12'd3566: q <= 1'b1;
			12'd3567: q <= 1'b1;
			12'd3568: q <= 1'b1;
			12'd3569: q <= 1'b1;
			12'd3570: q <= 1'b1;
			12'd3571: q <= 1'b1;
			12'd3572: q <= 1'b1;
			12'd3573: q <= 1'b1;
			12'd3574: q <= 1'b1;
			12'd3575: q <= 1'b1;
			12'd3576: q <= 1'b1;
			12'd3577: q <= 1'b0;
			12'd3578: q <= 1'b0;
			12'd3579: q <= 1'b0;
			12'd3580: q <= 1'b0;
			12'd3581: q <= 1'b0;
			12'd3582: q <= 1'b1;
			12'd3583: q <= 1'b1;
			12'd3584: q <= 1'b1;
			12'd3585: q <= 1'b1;
			12'd3586: q <= 1'b0;
			12'd3587: q <= 1'b1;
			12'd3588: q <= 1'b1;
			12'd3589: q <= 1'b1;
			12'd3590: q <= 1'b1;
			12'd3591: q <= 1'b1;
			12'd3592: q <= 1'b1;
			12'd3593: q <= 1'b1;
			12'd3594: q <= 1'b1;
			12'd3595: q <= 1'b1;
			12'd3596: q <= 1'b1;
			12'd3597: q <= 1'b1;
			12'd3598: q <= 1'b1;
			12'd3599: q <= 1'b1;
			12'd3600: q <= 1'b1;
			12'd3601: q <= 1'b1;
			12'd3602: q <= 1'b1;
			12'd3603: q <= 1'b1;
			12'd3604: q <= 1'b1;
			12'd3605: q <= 1'b1;
			12'd3606: q <= 1'b1;
			12'd3607: q <= 1'b1;
			12'd3608: q <= 1'b1;
			12'd3609: q <= 1'b1;
			12'd3610: q <= 1'b1;
			12'd3611: q <= 1'b1;
			12'd3612: q <= 1'b1;
			12'd3613: q <= 1'b1;
			12'd3614: q <= 1'b1;
			12'd3615: q <= 1'b1;
			12'd3616: q <= 1'b1;
			12'd3617: q <= 1'b0;
			12'd3618: q <= 1'b0;
			12'd3619: q <= 1'b0;
			12'd3620: q <= 1'b0;
			12'd3621: q <= 1'b0;
			12'd3622: q <= 1'b1;
			12'd3623: q <= 1'b1;
			12'd3624: q <= 1'b1;
			12'd3625: q <= 1'b1;
			12'd3626: q <= 1'b0;
			12'd3627: q <= 1'b1;
			12'd3628: q <= 1'b1;
			12'd3629: q <= 1'b1;
			12'd3630: q <= 1'b1;
			12'd3631: q <= 1'b1;
			12'd3632: q <= 1'b1;
			12'd3633: q <= 1'b1;
			12'd3634: q <= 1'b1;
			12'd3635: q <= 1'b1;
			12'd3636: q <= 1'b1;
			12'd3637: q <= 1'b1;
			12'd3638: q <= 1'b1;
			12'd3639: q <= 1'b1;
			12'd3640: q <= 1'b1;
			12'd3641: q <= 1'b1;
			12'd3642: q <= 1'b1;
			12'd3643: q <= 1'b1;
			12'd3644: q <= 1'b1;
			12'd3645: q <= 1'b1;
			12'd3646: q <= 1'b1;
			12'd3647: q <= 1'b1;
			12'd3648: q <= 1'b1;
			12'd3649: q <= 1'b1;
			12'd3650: q <= 1'b1;
			12'd3651: q <= 1'b1;
			12'd3652: q <= 1'b1;
			12'd3653: q <= 1'b1;
			12'd3654: q <= 1'b1;
			12'd3655: q <= 1'b1;
			12'd3656: q <= 1'b1;
			12'd3657: q <= 1'b0;
			12'd3658: q <= 1'b0;
			12'd3659: q <= 1'b0;
			12'd3660: q <= 1'b0;
			12'd3661: q <= 1'b0;
			12'd3662: q <= 1'b0;
			12'd3663: q <= 1'b1;
			12'd3664: q <= 1'b1;
			12'd3665: q <= 1'b1;
			12'd3666: q <= 1'b0;
			12'd3667: q <= 1'b1;
			12'd3668: q <= 1'b1;
			12'd3669: q <= 1'b1;
			12'd3670: q <= 1'b1;
			12'd3671: q <= 1'b1;
			12'd3672: q <= 1'b1;
			12'd3673: q <= 1'b1;
			12'd3674: q <= 1'b1;
			12'd3675: q <= 1'b1;
			12'd3676: q <= 1'b1;
			12'd3677: q <= 1'b1;
			12'd3678: q <= 1'b1;
			12'd3679: q <= 1'b1;
			12'd3680: q <= 1'b1;
			12'd3681: q <= 1'b1;
			12'd3682: q <= 1'b1;
			12'd3683: q <= 1'b1;
			12'd3684: q <= 1'b1;
			12'd3685: q <= 1'b1;
			12'd3686: q <= 1'b1;
			12'd3687: q <= 1'b1;
			12'd3688: q <= 1'b1;
			12'd3689: q <= 1'b1;
			12'd3690: q <= 1'b1;
			12'd3691: q <= 1'b1;
			12'd3692: q <= 1'b1;
			12'd3693: q <= 1'b1;
			12'd3694: q <= 1'b1;
			12'd3695: q <= 1'b1;
			12'd3696: q <= 1'b1;
			12'd3697: q <= 1'b0;
			12'd3698: q <= 1'b0;
			12'd3699: q <= 1'b0;
			12'd3700: q <= 1'b1;
			12'd3701: q <= 1'b1;
			12'd3702: q <= 1'b1;
			12'd3703: q <= 1'b1;
			12'd3704: q <= 1'b1;
			12'd3705: q <= 1'b1;
			12'd3706: q <= 1'b0;
			12'd3707: q <= 1'b1;
			12'd3708: q <= 1'b1;
			12'd3709: q <= 1'b1;
			12'd3710: q <= 1'b1;
			12'd3711: q <= 1'b1;
			12'd3712: q <= 1'b1;
			12'd3713: q <= 1'b1;
			12'd3714: q <= 1'b1;
			12'd3715: q <= 1'b1;
			12'd3716: q <= 1'b1;
			12'd3717: q <= 1'b1;
			12'd3718: q <= 1'b1;
			12'd3719: q <= 1'b1;
			12'd3720: q <= 1'b1;
			12'd3721: q <= 1'b1;
			12'd3722: q <= 1'b1;
			12'd3723: q <= 1'b1;
			12'd3724: q <= 1'b1;
			12'd3725: q <= 1'b1;
			12'd3726: q <= 1'b1;
			12'd3727: q <= 1'b1;
			12'd3728: q <= 1'b1;
			12'd3729: q <= 1'b1;
			12'd3730: q <= 1'b1;
			12'd3731: q <= 1'b1;
			12'd3732: q <= 1'b1;
			12'd3733: q <= 1'b1;
			12'd3734: q <= 1'b1;
			12'd3735: q <= 1'b1;
			12'd3736: q <= 1'b1;
			12'd3737: q <= 1'b0;
			12'd3738: q <= 1'b0;
			12'd3739: q <= 1'b0;
			12'd3740: q <= 1'b0;
			12'd3741: q <= 1'b0;
			12'd3742: q <= 1'b1;
			12'd3743: q <= 1'b1;
			12'd3744: q <= 1'b1;
			12'd3745: q <= 1'b1;
			12'd3746: q <= 1'b0;
			12'd3747: q <= 1'b1;
			12'd3748: q <= 1'b1;
			12'd3749: q <= 1'b1;
			12'd3750: q <= 1'b1;
			12'd3751: q <= 1'b1;
			12'd3752: q <= 1'b1;
			12'd3753: q <= 1'b1;
			12'd3754: q <= 1'b1;
			12'd3755: q <= 1'b1;
			12'd3756: q <= 1'b1;
			12'd3757: q <= 1'b1;
			12'd3758: q <= 1'b1;
			12'd3759: q <= 1'b1;
			12'd3760: q <= 1'b1;
			12'd3761: q <= 1'b1;
			12'd3762: q <= 1'b1;
			12'd3763: q <= 1'b1;
			12'd3764: q <= 1'b1;
			12'd3765: q <= 1'b1;
			12'd3766: q <= 1'b1;
			12'd3767: q <= 1'b1;
			12'd3768: q <= 1'b1;
			12'd3769: q <= 1'b1;
			12'd3770: q <= 1'b1;
			12'd3771: q <= 1'b1;
			12'd3772: q <= 1'b1;
			12'd3773: q <= 1'b1;
			12'd3774: q <= 1'b1;
			12'd3775: q <= 1'b1;
			12'd3776: q <= 1'b0;
			12'd3777: q <= 1'b0;
			12'd3778: q <= 1'b0;
			12'd3779: q <= 1'b0;
			12'd3780: q <= 1'b0;
			12'd3781: q <= 1'b0;
			12'd3782: q <= 1'b1;
			12'd3783: q <= 1'b1;
			12'd3784: q <= 1'b1;
			12'd3785: q <= 1'b1;
			12'd3786: q <= 1'b1;
			12'd3787: q <= 1'b1;
			12'd3788: q <= 1'b1;
			12'd3789: q <= 1'b1;
			12'd3790: q <= 1'b1;
			12'd3791: q <= 1'b1;
			12'd3792: q <= 1'b1;
			12'd3793: q <= 1'b1;
			12'd3794: q <= 1'b1;
			12'd3795: q <= 1'b1;
			12'd3796: q <= 1'b1;
			12'd3797: q <= 1'b1;
			12'd3798: q <= 1'b1;
			12'd3799: q <= 1'b1;
			12'd3800: q <= 1'b1;
			12'd3801: q <= 1'b1;
			12'd3802: q <= 1'b1;
			12'd3803: q <= 1'b1;
			12'd3804: q <= 1'b1;
			12'd3805: q <= 1'b1;
			12'd3806: q <= 1'b1;
			12'd3807: q <= 1'b1;
			12'd3808: q <= 1'b1;
			12'd3809: q <= 1'b1;
			12'd3810: q <= 1'b1;
			12'd3811: q <= 1'b1;
			12'd3812: q <= 1'b1;
			12'd3813: q <= 1'b1;
			12'd3814: q <= 1'b1;
			12'd3815: q <= 1'b1;
			12'd3816: q <= 1'b0;
			12'd3817: q <= 1'b0;
			12'd3818: q <= 1'b0;
			12'd3819: q <= 1'b0;
			12'd3820: q <= 1'b0;
			12'd3821: q <= 1'b0;
			12'd3822: q <= 1'b0;
			12'd3823: q <= 1'b1;
			12'd3824: q <= 1'b1;
			12'd3825: q <= 1'b1;
			12'd3826: q <= 1'b1;
			12'd3827: q <= 1'b0;
			12'd3828: q <= 1'b1;
			12'd3829: q <= 1'b1;
			12'd3830: q <= 1'b1;
			12'd3831: q <= 1'b1;
			12'd3832: q <= 1'b1;
			12'd3833: q <= 1'b1;
			12'd3834: q <= 1'b1;
			12'd3835: q <= 1'b1;
			12'd3836: q <= 1'b1;
			12'd3837: q <= 1'b1;
			12'd3838: q <= 1'b1;
			12'd3839: q <= 1'b1;
			12'd3840: q <= 1'b1;
			12'd3841: q <= 1'b1;
			12'd3842: q <= 1'b1;
			12'd3843: q <= 1'b1;
			12'd3844: q <= 1'b1;
			12'd3845: q <= 1'b1;
			12'd3846: q <= 1'b1;
			12'd3847: q <= 1'b1;
			12'd3848: q <= 1'b1;
			12'd3849: q <= 1'b1;
			12'd3850: q <= 1'b1;
			12'd3851: q <= 1'b1;
			12'd3852: q <= 1'b1;
			12'd3853: q <= 1'b1;
			12'd3854: q <= 1'b1;
			12'd3855: q <= 1'b0;
			12'd3856: q <= 1'b0;
			12'd3857: q <= 1'b0;
			12'd3858: q <= 1'b0;
			12'd3859: q <= 1'b0;
			12'd3860: q <= 1'b0;
			12'd3861: q <= 1'b0;
			12'd3862: q <= 1'b0;
			12'd3863: q <= 1'b1;
			12'd3864: q <= 1'b1;
			12'd3865: q <= 1'b1;
			12'd3866: q <= 1'b1;
			12'd3867: q <= 1'b1;
			12'd3868: q <= 1'b1;
			12'd3869: q <= 1'b0;
			12'd3870: q <= 1'b0;
			12'd3871: q <= 1'b1;
			12'd3872: q <= 1'b1;
			12'd3873: q <= 1'b1;
			12'd3874: q <= 1'b1;
			12'd3875: q <= 1'b1;
			12'd3876: q <= 1'b1;
			12'd3877: q <= 1'b1;
			12'd3878: q <= 1'b1;
			12'd3879: q <= 1'b1;
			12'd3880: q <= 1'b1;
			12'd3881: q <= 1'b1;
			12'd3882: q <= 1'b1;
			12'd3883: q <= 1'b1;
			12'd3884: q <= 1'b1;
			12'd3885: q <= 1'b1;
			12'd3886: q <= 1'b1;
			12'd3887: q <= 1'b1;
			12'd3888: q <= 1'b1;
			12'd3889: q <= 1'b1;
			12'd3890: q <= 1'b1;
			12'd3891: q <= 1'b1;
			12'd3892: q <= 1'b0;
			12'd3893: q <= 1'b0;
			12'd3894: q <= 1'b0;
			12'd3895: q <= 1'b0;
			12'd3896: q <= 1'b0;
			12'd3897: q <= 1'b0;
			12'd3898: q <= 1'b0;
			12'd3899: q <= 1'b0;
			12'd3900: q <= 1'b0;
			12'd3901: q <= 1'b0;
			12'd3902: q <= 1'b0;
			12'd3903: q <= 1'b1;
			12'd3904: q <= 1'b1;
			12'd3905: q <= 1'b0;
			12'd3906: q <= 1'b0;
			12'd3907: q <= 1'b0;
			12'd3908: q <= 1'b0;
			12'd3909: q <= 1'b0;
			12'd3910: q <= 1'b0;
			12'd3911: q <= 1'b0;
			12'd3912: q <= 1'b0;
			12'd3913: q <= 1'b0;
			12'd3914: q <= 1'b0;
			12'd3915: q <= 1'b1;
			12'd3916: q <= 1'b1;
			12'd3917: q <= 1'b1;
			12'd3918: q <= 1'b1;
			12'd3919: q <= 1'b1;
			12'd3920: q <= 1'b0;
			12'd3921: q <= 1'b0;
			12'd3922: q <= 1'b0;
			12'd3923: q <= 1'b0;
			12'd3924: q <= 1'b0;
			12'd3925: q <= 1'b0;
			12'd3926: q <= 1'b0;
			12'd3927: q <= 1'b0;
			12'd3928: q <= 1'b0;
			12'd3929: q <= 1'b0;
			12'd3930: q <= 1'b0;
			12'd3931: q <= 1'b0;
			12'd3932: q <= 1'b0;
			12'd3933: q <= 1'b0;
			12'd3934: q <= 1'b0;
			12'd3935: q <= 1'b0;
			12'd3936: q <= 1'b0;
			12'd3937: q <= 1'b0;
			12'd3938: q <= 1'b0;
			12'd3939: q <= 1'b0;
			12'd3940: q <= 1'b0;
			12'd3941: q <= 1'b0;
			12'd3942: q <= 1'b0;
			12'd3943: q <= 1'b0;
			12'd3944: q <= 1'b0;
			12'd3945: q <= 1'b0;
			12'd3946: q <= 1'b0;
			12'd3947: q <= 1'b0;
			12'd3948: q <= 1'b0;
			12'd3949: q <= 1'b0;
			12'd3950: q <= 1'b0;
			12'd3951: q <= 1'b0;
			12'd3952: q <= 1'b0;
			12'd3953: q <= 1'b0;
			12'd3954: q <= 1'b0;
			12'd3955: q <= 1'b0;
			12'd3956: q <= 1'b0;
			12'd3957: q <= 1'b0;
			12'd3958: q <= 1'b0;
			12'd3959: q <= 1'b0;
			12'd3960: q <= 1'b0;
			12'd3961: q <= 1'b0;
			12'd3962: q <= 1'b0;
			12'd3963: q <= 1'b0;
			12'd3964: q <= 1'b0;
			12'd3965: q <= 1'b0;
			12'd3966: q <= 1'b0;
			12'd3967: q <= 1'b0;
			12'd3968: q <= 1'b0;
			12'd3969: q <= 1'b0;
			12'd3970: q <= 1'b0;
			12'd3971: q <= 1'b0;
			12'd3972: q <= 1'b0;
			12'd3973: q <= 1'b0;
			12'd3974: q <= 1'b0;
			12'd3975: q <= 1'b0;
			12'd3976: q <= 1'b0;
			12'd3977: q <= 1'b0;
			12'd3978: q <= 1'b0;
			12'd3979: q <= 1'b0;
			12'd3980: q <= 1'b0;
			12'd3981: q <= 1'b0;
			12'd3982: q <= 1'b0;
			12'd3983: q <= 1'b0;
			12'd3984: q <= 1'b0;
			12'd3985: q <= 1'b0;
			12'd3986: q <= 1'b0;
			12'd3987: q <= 1'b0;
			12'd3988: q <= 1'b0;
			12'd3989: q <= 1'b0;
			12'd3990: q <= 1'b0;
			12'd3991: q <= 1'b0;
			12'd3992: q <= 1'b0;
			12'd3993: q <= 1'b0;
			12'd3994: q <= 1'b0;
			12'd3995: q <= 1'b0;
			12'd3996: q <= 1'b1;
			12'd3997: q <= 1'b1;
			12'd3998: q <= 1'b1;
			12'd3999: q <= 1'b1;
		endcase	
	end
	assign out = q;
endmodule