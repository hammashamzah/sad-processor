module without_uart_testbench();

	reg clk;
	reg rst;
	reg UARTstart;
	reg UARTready;
	reg UARTsendComplete;
	reg[7:0] data_in;
	
	wire valid;
	wire[9:0] x_out;
	wire[8:0] y_out;
	wire[7:0] data_in_reverse;

	topLevel_withoutUART toplevel
	(
		.clock(clk),
		.reset(rst),
		.UARTstart(UARTstart),
		.UARTready(UARTready),
		.UARTsendComplete(UARTsendComplete),
		.data_in(data_in_reverse),
		.valid(valid),
		.x_out(x_out),
		.y_out(y_out)
	);
	
	genvar i;
	generate
		for (i = 0; i < 8; i = i + 1)
		begin:reverse
			assign data_in_reverse[i] = data_in[7 - i];			
		end
	endgenerate


	/** Clock generation **/
	always
		#5 clk = ~clk;
	
	/** Send inputs and receive outputs **/
	initial
	begin
		clk   = 1'b1;
		rst   = 1'b1;
		UARTsendComplete = 1'b0;
		UARTstart = 1'b0;
		UARTready = 1'b0;
		#20
		rst = 1'b0;
		#10
		UARTstart = 1'b1;
		#10
		UARTstart = 1'b0;
		
		#10
		UARTready = 1'b1;

		data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b00010001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10010000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b10010011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b11011111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b10000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10001011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b11000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01010111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b11101111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010111;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b01011011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00100011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01101111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11110110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01101111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11001110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11101111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11101111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11011110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11011110;
		#10 data_in[7:0] =  8'b01111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b01111100;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b01001100;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111010;
		#10 data_in[7:0] =  8'b00111100;
		#10 data_in[7:0] =  8'b10011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b01001000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111010;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b01111010;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01110000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01110001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01110110;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01110000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01110000;
		#10 data_in[7:0] =  8'b01110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b10011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b01100110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b00001001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001011;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001011;
		#10 data_in[7:0] =  8'b01110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11100011;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111011;
		#10 data_in[7:0] =  8'b11011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11011011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100011;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01110000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01100011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b10101111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11011001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110001;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11100011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b11011001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10111000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11001001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100010;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11001011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11101111;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11001001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10011000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b10111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01100011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111010;
		#10 data_in[7:0] =  8'b11000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b10111100;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b00110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110110;
		#10 data_in[7:0] =  8'b01010011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10011000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10011000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b00010011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10011111;
		#10 data_in[7:0] =  8'b01100001;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01101111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10001100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b10010011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10010100;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b10011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111110;
		#10 data_in[7:0] =  8'b00011100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11010011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11110100;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00011100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000101;
		#10 data_in[7:0] =  8'b11111001;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11010011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b10000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11001101;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10111110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11010011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b10001100;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10010011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b01111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b01001110;
		#10 data_in[7:0] =  8'b01110000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11010011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00101111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11011110;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00111011;
		#10 data_in[7:0] =  8'b11000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b11001100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100001;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b11001110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010010;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b11000110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b10000010;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000101;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b10010011;
		#10 data_in[7:0] =  8'b11110110;
		#10 data_in[7:0] =  8'b10010101;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b01111101;
		#10 data_in[7:0] =  8'b11000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b10000010;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11000100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10010011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11001001;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00111101;
		#10 data_in[7:0] =  8'b11000011;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000010;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01010011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111001;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00111101;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000110;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b10100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11011011;
		#10 data_in[7:0] =  8'b11000111;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b10111001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000101;
		#10 data_in[7:0] =  8'b11101111;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b10000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00111001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00001110;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b10000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b10111001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11110001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b10101110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111011;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b01111110;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010011;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110011;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110011;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00101100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111110;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11110001;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11101101;
		#10 data_in[7:0] =  8'b10011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b01111011;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00011100;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00001110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b01001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00001110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00001110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00001110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000101;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b10000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011100;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100010;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b10000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010110;
		#10 data_in[7:0] =  8'b01100100;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01001111;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01011110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11000101;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b10000111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00011100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01011110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11011111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b00011100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00010011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01011110;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b10011111;
		#10 data_in[7:0] =  8'b11010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10001000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b01110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011101;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b01110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11000011;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b01110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00111011;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001011;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11000011;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000110;
		#10 data_in[7:0] =  8'b10001100;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10100111;
		#10 data_in[7:0] =  8'b10000101;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100001;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b01110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000111;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b10001100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100001;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100011;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100001;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b10100001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b10001111;
		#10 data_in[7:0] =  8'b01110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000101;
		#10 data_in[7:0] =  8'b10000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100011;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10111100;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b01111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110110;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b10000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b01111110;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01001111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011011;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001011;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000111;
		#10 data_in[7:0] =  8'b11011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00001110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111010;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00111010;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00001110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00001110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b01111101;
		#10 data_in[7:0] =  8'b10100110;
		#10 data_in[7:0] =  8'b11000010;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11101100;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11101000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b10000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00011100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111010;
		#10 data_in[7:0] =  8'b01111000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11101111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b01111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b11000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00011100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111010;
		#10 data_in[7:0] =  8'b01111100;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b00111010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111010;
		#10 data_in[7:0] =  8'b11110100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11101100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00011000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b01111010;
		#10 data_in[7:0] =  8'b00111100;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b10111000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b10111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00011000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111000;
		#10 data_in[7:0] =  8'b00111000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11101000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b00001101;
		#10 data_in[7:0] =  8'b11100100;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11101111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00100100;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100011;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11011000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10011100;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01011111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00111001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b11000111;
		#10 data_in[7:0] =  8'b10110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011100;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b10011111;
		#10 data_in[7:0] =  8'b01001111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110100;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00011001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b01011010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00001001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b00001011;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b00100111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00011011;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01110000;
		#10 data_in[7:0] =  8'b00011000;
		#10 data_in[7:0] =  8'b00011001;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b10000111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100001;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b00111100;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111011;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001011;
		#10 data_in[7:0] =  8'b00001101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10100101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11101000;
		#10 data_in[7:0] =  8'b01111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b01111100;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b00010111;
		#10 data_in[7:0] =  8'b00010111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11000001;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01011111;
		#10 data_in[7:0] =  8'b11010110;
		#10 data_in[7:0] =  8'b10000011;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00111110;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111110;
		#10 data_in[7:0] =  8'b00001110;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11110001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00101111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000101;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b01000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00001011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010100;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11101111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01110000;
		#10 data_in[7:0] =  8'b00010011;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10101011;
		#10 data_in[7:0] =  8'b11001000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b01110111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b11110001;
		#10 data_in[7:0] =  8'b11000001;
		#10 data_in[7:0] =  8'b00101000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000001;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11100011;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00101111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011010;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00101111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00011000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00011100;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11001000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11101101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b00000101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b10110111;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011100;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10010000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11011000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b00000101;
		#10 data_in[7:0] =  8'b01101111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01011000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b01111101;
		#10 data_in[7:0] =  8'b01111110;
		#10 data_in[7:0] =  8'b11011001;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b10011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00011100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001011;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b01110000;
		#10 data_in[7:0] =  8'b01000010;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10011000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11101000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00011011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100011;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b10000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01101100;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b10010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01110100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001001;
		#10 data_in[7:0] =  8'b10000011;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b10001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b01101100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01001110;
		#10 data_in[7:0] =  8'b11000001;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b01011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11101110;
		#10 data_in[7:0] =  8'b00100001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b00101110;
		#10 data_in[7:0] =  8'b11000011;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000011;
		#10 data_in[7:0] =  8'b10111110;
		#10 data_in[7:0] =  8'b00010100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11000011;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b01111101;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b01111110;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b10011000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001110;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11110110;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b10100000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11000011;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000011;
		#10 data_in[7:0] =  8'b10010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11011110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111110;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11001000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000011;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10011111;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111001;
		#10 data_in[7:0] =  8'b01111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000011;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b01011111;
		#10 data_in[7:0] =  8'b11010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b00111100;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111110;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00011000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000011;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b01001111;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00011100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010110;
		#10 data_in[7:0] =  8'b00100111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b01111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01001111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01010111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100001;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b10001000;
		#10 data_in[7:0] =  8'b01101000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10110001;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110110;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111110;
		#10 data_in[7:0] =  8'b01111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11101111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000110;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11000001;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00110010;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11101111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b11100001;
		#10 data_in[7:0] =  8'b11110110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000011;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b11001100;
		#10 data_in[7:0] =  8'b00000101;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01100001;
		#10 data_in[7:0] =  8'b01111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b10000011;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b10011111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000111;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11000001;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110110;
		#10 data_in[7:0] =  8'b01101110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b01011100;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111001;
		#10 data_in[7:0] =  8'b00111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00101111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100001;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00010001;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b10000101;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11010111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00001110;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11110100;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11011111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10010110;
		#10 data_in[7:0] =  8'b00010001;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11101111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001110;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000011;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11100011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b10100000;
		#10 data_in[7:0] =  8'b00011000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00011000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b01111110;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b10011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11001110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b10010001;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01011110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011011;
		#10 data_in[7:0] =  8'b11010000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b10110001;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100011;
		#10 data_in[7:0] =  8'b10111101;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b10110000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110011;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11000100;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b01111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011101;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b10000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110111;
		#10 data_in[7:0] =  8'b00111101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111000;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000101;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b00001110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11110001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b11000100;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11110001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111000;
		#10 data_in[7:0] =  8'b00011000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111100;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11110110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11100010;
		#10 data_in[7:0] =  8'b00011000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11101100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b11011000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11101111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b01111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00001011;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01110111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b11100100;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10011100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b10000111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00101000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011100;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11100011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b10001000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111110;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10101111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11000010;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11101011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b10011000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11001100;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b01001001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b01001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11011110;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00111011;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b10100000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01110000;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11101000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111100;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b01111110;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b11101100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111110;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b10000011;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010001;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00101111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01011110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111011;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b11101111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00011000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01110010;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b01101000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b00001010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00011000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10011101;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111000;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111110;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b01100111;
		#10 data_in[7:0] =  8'b11110110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011101;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b10000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00011000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b10100000;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00001011;
		#10 data_in[7:0] =  8'b01010110;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01110011;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01110000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b11111001;
		#10 data_in[7:0] =  8'b11110100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b11000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01110000;
		#10 data_in[7:0] =  8'b01111110;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b01011101;
		#10 data_in[7:0] =  8'b10000110;
		#10 data_in[7:0] =  8'b00001001;
		#10 data_in[7:0] =  8'b11100001;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b11011111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b10000110;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b01011100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10101111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b10011111;
		#10 data_in[7:0] =  8'b11000011;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000001;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11100011;
		#10 data_in[7:0] =  8'b10111011;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00010011;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000001;
		#10 data_in[7:0] =  8'b00111110;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b11011110;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01110000;
		#10 data_in[7:0] =  8'b00100111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10001000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11100011;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11011111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b01111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111010;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b11000001;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11101101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11001000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b01110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11011000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00011000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001110;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100111;
		#10 data_in[7:0] =  8'b10111110;
		#10 data_in[7:0] =  8'b01100111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b01000111;
		#10 data_in[7:0] =  8'b10111110;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b10111000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b10011111;
		#10 data_in[7:0] =  8'b10111110;
		#10 data_in[7:0] =  8'b00101111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b10011111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b11110001;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b10001111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111001;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00100001;
		#10 data_in[7:0] =  8'b11011111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01011111;
		#10 data_in[7:0] =  8'b11010000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00010100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b10100000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11110001;
		#10 data_in[7:0] =  8'b11010101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111101;
		#10 data_in[7:0] =  8'b11110101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b11100110;
		#10 data_in[7:0] =  8'b01111001;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11011111;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b01000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10011111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100111;
		#10 data_in[7:0] =  8'b11101111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111000;
		#10 data_in[7:0] =  8'b10010001;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00100111;
		#10 data_in[7:0] =  8'b10001111;
		#10 data_in[7:0] =  8'b11111001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b10011111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11101111;
		#10 data_in[7:0] =  8'b10110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11100110;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b10000110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11100010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00101111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11101011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00010110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01100001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111010;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010110;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000100;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00110010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b00011001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b01110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b01110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b01111000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b10111011;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11000111;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b01011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b01001000;
		#10 data_in[7:0] =  8'b11000111;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00101111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001110;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011011;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11001011;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10011111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00001110;
		#10 data_in[7:0] =  8'b11011111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b11000011;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10001111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b10001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000101;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000101;
		#10 data_in[7:0] =  8'b10100111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11001011;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b01111100;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11100001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10011111;
		#10 data_in[7:0] =  8'b01110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11100011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00001110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11101111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b10000011;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00111101;
		#10 data_in[7:0] =  8'b10000111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00001101;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b11010000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11001100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111100;
		#10 data_in[7:0] =  8'b00001110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11110100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b00001110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10001111;
		#10 data_in[7:0] =  8'b11100101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000001;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b01100111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10100100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b01111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100011;
		#10 data_in[7:0] =  8'b00011000;
		#10 data_in[7:0] =  8'b00101111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b01111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11000110;
		#10 data_in[7:0] =  8'b00011010;
		#10 data_in[7:0] =  8'b01110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b01111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11011111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b01111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011101;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111010;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b01011111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b00111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00100011;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b01100100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11110101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000001;
		#10 data_in[7:0] =  8'b01000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01011100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b00011000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b10001001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b00100110;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111000;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11000110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00101000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01100110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01110001;
		#10 data_in[7:0] =  8'b11011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b01111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00001110;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b00101111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b01110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11000001;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11011110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b11101100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11011111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10001100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11101111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b00010111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110001;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00001110;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111001;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b01111100;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00111110;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11101111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b10011100;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b10111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11010000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001110;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b11101111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011100;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11101111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11100001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111010;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00110100;
		#10 data_in[7:0] =  8'b11101111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100001;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111100;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00111100;
		#10 data_in[7:0] =  8'b01101111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000101;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b01110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b10011110;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11100010;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b01011100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11011110;
		#10 data_in[7:0] =  8'b10100000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10011110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000010;
		#10 data_in[7:0] =  8'b01101000;
		#10 data_in[7:0] =  8'b11001101;
		#10 data_in[7:0] =  8'b11110001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00111110;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00001110;
		#10 data_in[7:0] =  8'b01100111;
		#10 data_in[7:0] =  8'b10001001;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10111110;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00001010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11000001;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b00001001;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111100;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000110;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011110;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11000011;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011100;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b10011111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010010;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01110000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001101;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11100001;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11010000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b10000111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110011;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10010101;
		#10 data_in[7:0] =  8'b10000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011100;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001110;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111010;
		#10 data_in[7:0] =  8'b10000011;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b11000011;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001001;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b11101100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11101111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11101111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11101001;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10011111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111010;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11101111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b10110001;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111100;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b01110011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111101;
		#10 data_in[7:0] =  8'b11101000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011100;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b11000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11100001;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111000;
		#10 data_in[7:0] =  8'b01010000;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10100000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11001000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11101111;
		#10 data_in[7:0] =  8'b11011000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b10000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b11111010;
		#10 data_in[7:0] =  8'b10011111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10010111;
		#10 data_in[7:0] =  8'b00001011;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01110000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11110001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000010;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111011;
		#10 data_in[7:0] =  8'b01000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00011010;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110111;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00110011;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b11011111;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11101000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11001000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b10011100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111101;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01101000;
		#10 data_in[7:0] =  8'b00001100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01100011;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b10111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b10100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000110;
		#10 data_in[7:0] =  8'b01110011;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b10011111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b00011001;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01100001;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11000001;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00011000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11110001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010011;
		#10 data_in[7:0] =  8'b11111101;
		#10 data_in[7:0] =  8'b11011111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b10110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b01000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00010111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10100100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11101000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111110;
		#10 data_in[7:0] =  8'b01100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b01110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000001;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111010;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111100;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11001111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b10000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00001000;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11101111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11100000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000100;
		#10 data_in[7:0] =  8'b00111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b01111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000011;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11110000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00000000;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b00011111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 data_in[7:0] =  8'b11111111;
		#10 UARTready = 1'b0;


	end
	
endmodule 