module original_image_rom(
	input	[8:0]addr,
	input	clk,
	output	[639:0]out
);
	reg [639:0]q;

	always @(posedge clk)
	begin
		case(addr)
			9'd 00: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 01: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 02: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 03: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 04: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 05: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 06: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 07: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 08: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 09: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 10: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 11: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 12: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 13: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 14: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 15: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 16: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 17: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 18: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 19: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 20: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 21: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 22: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 23: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 24: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 25: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 26: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 27: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 28: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 29: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 30: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 31: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 32: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 33: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 34: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 35: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 36: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 37: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 38: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 39: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 40: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 41: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 42: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 43: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 44: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 45: q <= 640'b1111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 46: q <= 640'b1111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 47: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 48: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 49: q <= 640'b1111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 50: q <= 640'b1111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 51: q <= 640'b1111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 52: q <= 640'b1111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 53: q <= 640'b1111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 54: q <= 640'b1111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 55: q <= 640'b1111111111111111111011111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 56: q <= 640'b1111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 57: q <= 640'b1111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 58: q <= 640'b1111111111111111111001111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 59: q <= 640'b1111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 60: q <= 640'b1111111111111111111000000000100111111111100010001100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 61: q <= 640'b1111111111111111111000000000000111111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 62: q <= 640'b1111111111111111111000000000000011111000001111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 63: q <= 640'b1111111111111111111001111111111111110000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 64: q <= 640'b1111111111111111111001111111111111111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 65: q <= 640'b1111111111111111111001111111111111111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 66: q <= 640'b1111111111111111110001111111111111111000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 67: q <= 640'b1111111111111111111001111111111111111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 68: q <= 640'b1111111111111111111001111111111111111011111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 69: q <= 640'b1111111111111111101001111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 70: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 71: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 72: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 73: q <= 640'b1111111111111111111111110011111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 74: q <= 640'b1111101111111111110010010011111111111101000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 75: q <= 640'b1111101111111111110000010011111111111011000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 76: q <= 640'b1111111111111111111000110001111111111110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 77: q <= 640'b1111111111111111111101110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 78: q <= 640'b0111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 79: q <= 640'b0110111111111111111110010000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 80: q <= 640'b1110100000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 81: q <= 640'b1111110111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111;
			9'd 82: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 83: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 84: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 85: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 86: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 87: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000100000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 88: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 89: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 90: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 91: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 92: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 93: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 94: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 95: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 96: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 97: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 98: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd 99: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd100: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd101: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111111111111000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd102: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd103: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd104: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101111111111000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
			9'd105: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000111111111100001111111111111111111111111111111111111111111111111111111111111111111111;
			9'd106: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110011111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000001111110000000011111111111111111111111111111111111111111111111111111111111111111111;
			9'd107: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111001110000000011111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111000000000001111111111111111111111111111111111111111111111111111111111111111111;
			9'd108: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111011111111111100000000011111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111110000000000001111111111111111111111111111111111111111111111111111111111111111111;
			9'd109: q <= 640'b1111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110011110110000000000011111111111111111111111111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000111110000000000000111111111111111111111111111111111111111111111111111111111111111111;
			9'd110: q <= 640'b1111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100001111100100000000111111111111111111111111111111111111111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000001111100000000000001111111111111111111111111111111111111111111111111111111111111111111;
			9'd111: q <= 640'b1111111111111001001111000101111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111001100110010000111111000000000011111111111111111111111111111111111111111111111111111111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000001111100000000000001111111111111111111111111111111111111111111111111111111111111111111;
			9'd112: q <= 640'b1111111111110011111111100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000010010000011111000000000000011111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000001111100000000000001111111111111111111111111111111111111111111111111111111111111111111;
			9'd113: q <= 640'b1111111111111111111111110101111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111000000000000000000010000001111110000000000001111111111111111111111111111111111111111111111111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000001111100000000000000111111111111111111111111111111111111111111111111111111111111100101;
			9'd114: q <= 640'b1111111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000111110110111000000000000000000000000000000000000011111111111111111111111111111111111111111111111111110000000000000000000000000000000000000010000000001000111000000000011111111111111111111111111111111111111111111111111111111111100000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000111000000000000000111111111111111111111111111111111111111111111111111111111111111111;
			9'd115: q <= 640'b1111111111111111100111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111110000000000000000000000000010000000000000000000000000000000010000010000000111000000000001111111111111111111111111111111111111111111111111111111111100000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111110;
			9'd116: q <= 640'b1111111111111111111100000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000000000000000000010000000000111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000111000001110000000000000000000000010000000000000110000000000001111111111111111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000111111111111111111111111111111111111111111111111111111111111001100;
			9'd117: q <= 640'b1111111111111111110000000000000000000011111110000000011111111111111111111111111111111111011001100111111111110011101111111111111111111111111111111111110000000000011111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000001111100011111000000000000000000000011000000000000000000000000000111111111111111111111111111111111111111111111111111111111000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000111111111111111001000001111000000000000000000000000000000000000000;
			9'd118: q <= 640'b1111111111111111110000000000000000000011111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111100000000000000000000011100000000000000000000000000111111111111111111111111111111111111111111111111111111111000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd119: q <= 640'b1111111111111111110000000000000000000011111100000000000111111111111111111101111111111111111111111111111111111111111111111111111111111111111111011101000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000000000011100000000000000000000000000111111111111111111111111111111111111111111111111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd120: q <= 640'b1111111111111111000000000000000000000011111000000000000111111111111111111101111111111111111111111111111111111110111100000000000000000000000011101101000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111100000000000000000000011100000000000000000000000000111111111111111111111111111111111111111111111111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd121: q <= 640'b1111111111101111000000000000000000000011111000000000000111111111111111111100001111111111111111101111111111111111111111111111111111111111111111111101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111100000000000000000000011100000000000000000000000000011111111111111111111111111111111111111111111111111111100000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111001100011111111100;
			9'd122: q <= 640'b1111111111110010000000000000000000000001111000000000000011111111111111111100111111111111111111111111111111111111111111111111111111111111111111111001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111100000000000000000000011100000000000000000000000110011111111111111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111011111111111111111111111111111111111111111111111111111;
			9'd123: q <= 640'b1111111111100100000000000000000000000101100000000000000011111111111111111101101111111111111111111100111111111111111111111111111111111111111110111101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111100000000000000000000011110000000000000000000000010111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111110000000000000001011110000000000000000000000000001111111111011111111111111111111111111111111111111111111111111111;
			9'd124: q <= 640'b1111111111100100000000000000000000000000001000000000000111111111111111111001101111111111111111111111000011111111111111111111010110111111111111111100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111110000000000000000000000011100000000000000000000000011011111111111111111111111111111111100000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000001111110001111111111111111111111111110000001111111111111111111100000000000000000000011111111111011111111111111111111111111111111111111111111111111111;
			9'd125: q <= 640'b1111111111111000000000000000000000000000000100000000000011111111111111111001101110111111111111111110000001111111111111111111110111111111111111111100011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111110000000000000000000000011110000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001111111100011111111111111111111111111111111111111111111111001111111111111111111111111110000001111111111111111111100000000000000000000011111111111011111111111111111111111111111111111111111111111111111;
			9'd126: q <= 640'b1111111111110000000000000000000000000000000100000000000001111111111111111001001111111111111111111100000000001111111111111101111111100111111111100001110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100011111110000000000000000000000011110000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111001111111111111111111111111110000001111111111111111111100000000000000000000011111111111111111111111111111111111111111111111111111111111111111;
			9'd127: q <= 640'b1111110010000000000000000000000000000000000010000000000011111111111111111101001111111111111111111100000000000011010001111111111111111111111111000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000011110000000000000000000001100000000000000000000000000000001111111011111111111111111100000000000000000001111111111111111111111111111111111111111111110011111111111111111111101111111111111111111111111001111111111111111111111111110000001111111111111111111100000000000000000000011111111110111111111111111111111111111111111111111111111111111111;
			9'd128: q <= 640'b1111101100000000000000000000000000000000000000000000000101111111111111111001001111111111111111111000000000000000000111111111110011110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000011000000000000000000000001001111111111111111111111111111101111111111111111111111111100000000000000000000111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111001111111111111111111111111110000001111111111111111111100000000000000000000111111111110011111111111111111111111111110111111111111111111111111;
			9'd129: q <= 640'b1110110010000000000000000000000000000000000001000000000111111111111111111100001101011111111111111100011000000000000011111111111111011101111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000011001000000000000000000000010011111111111111111111111111111101111111111111111111111111100000000000000000000011111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111001111111111111111111111111110000001111111111111111111100000000000000000000111111111110011111111111111111111111111111111111111111111111111111;
			9'd130: q <= 640'b1111100010000000000000000000000000000000000001100000001111111101111111111100101001101111111111111110110001100000000011111111111100111101111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000001000000000000000000000101111111111111111111111111111111101111111111111111111111111100000000000000000000001111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111001111111111111111111111111110000001111111111111111111110000000000000000000111111111110011111111111111111111111111111111111111111111111111111;
			9'd131: q <= 640'b1111011000000000000000000000000000000000000111111000011011111001111111111100100011101111111111111111101000000000000001111111111100011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000001000000000000000000011001111111111111111111111111111111101111111111111111111111111100000000000000000000000111111111111111111111111111111111111111110011111111111111111111101111111111111111111111111001111111111111111111111111110000011111111111111111111110000000000000000000111111111110011111111111111111111111111111111111111111111111111111;
			9'd132: q <= 640'b1111111000000000000000000000000000000000011111111111001111111111111111111100100111011111111111111101110000000010110111111111111100000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000001100000000000000000110001111111111111111111111111111111101111111111111111111111111000000000000000000000000111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111001111111111111111111111111110000011111111111111111111100000000000000000001111111111110011111111111111111111111111111111111111111111111111110;
			9'd133: q <= 640'b1111111000000000000000000000000000000001111111111111111011111101111111111100000011111111111111111111100111100000111111111111111000101001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000011111110000000000000000000000001100000000000000000100000111111111111111111111111111111101111111111111111111111110000000000000000000000000011111111111111111111111111111111111111110011111111111111111111111111111111111111111111111001111111111111111111111111110000011111111111111111111100000000000000000001111111111110011111111111111111111111111111111111111111111111111000;
			9'd134: q <= 640'b0010111100000000000000000000000000000011111111111111111111111111111111111100101111111111111111111111111111111100001111111111100000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001111110000000000000000000000001000000000000000000000000111111111111111111111111111111101111111111111111111111100000000000000000000000000001111111111111111111111111111111111111110011111111111111111111111111111111111111111111111011111111111111111111111111110000011111111111111111000000000000000000000011111111111110001111111111111111111111111111111111111111111111100000;
			9'd135: q <= 640'b1110000000000000000000000000000000000011111111111111111101111111111111111100101111111111111111111111111111101111100111111010000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001111111000000000000000000000001000000000000000000000000111111111111111111111111111111101111111111111111111111100000000000000000000000000000111111111111111111111111111111111111110011111111111111111111101111111111111111111111110011111111111111111111111111111000011111111111111100000000000000000000000011111111111110011111111111111111111111111111111111111111111110000000;
			9'd136: q <= 640'b1011001100000000000000000000000000000111111111111111111111111111111111111100001111111111111011111111111111100001111111010010000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000111111000000000000000000000001100000000000000000000000111111111111111111111111111111101111111111111111111111000000000000000000000000000000111111111111111111111111111111111111110011111111111111111111111111111111111111111111111011111111111111111111111111110000011111111000000000000000000000000000000011111111111110011111111111111111111111111111111111111111111000000000;
			9'd137: q <= 640'b0010100000000000000000000000000000001111111111111111111111111111111111111100101111111111111111111111111111111111011111011000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110001111111000000000000000000000001100000000000000000000000111111111111111111111111111111101111111111111111111110000000000000000000000000000000111111111111111111111111111111111111110011111111111111111111111111111111111111111111110011111111111111111111111111110000011111111111110000001000000000000000000011111111111100111111111111111111111111111111111111111111111000000000;
			9'd138: q <= 640'b1111110000000000000000000000000000011111111111111111111111111111111111111100100111111111111111111111111111111111001100011100000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000001111000000000000000000000001100000000000000000000000111111111111111111111111111111101111111111111111111100000000000000000000000000000000111111111111111111111111111111111111110011111111111111111111111111111111111111111111110011111111111111111111111111110000011111111111111100111000000000000000000001111111111100111111111111111111111111111111111111111111100000000000;
			9'd139: q <= 640'b1111111000000000000000000000000000111111111111111111101111111111111111111100101111111111111111111111111000001110011100101111100000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111001111000000000000000000000000001100000000000000000000000111111111111111111111111111111101111111101111111111100000000000000000000000000000000111111111111111111111111111111111111110011111111111111111111111111111111111111111111110011111111111111111111111111110000011111111111111111110000000000000000000011111111111100111111111111111111111111111111111111111111100000000000;
			9'd140: q <= 640'b1111100000000000000000000000000000110011101111111111001111111111111111111100111111111111111000111101110000000011011110111111100000000111001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000000000000111111111111111111111111111111111111111111111111111101000000000000000000000000000000011111111111111111111111111111111111110011111111111111111111111111111111111111111111110011111111111111111111111111110000011111111111111111100000000000000000000011111111111000011111111111111111111111111111111111111111000000000000;
			9'd141: q <= 640'b1111111000000000000000000000000001110011101111111000011111111111111111111100100000000000000001111111110000000000001111111111100000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000100000000000001111111111111111111111111111111111111111111111111111111000000000000000000000000000000011111111111111111111111111111111111110011111111111111111111111111111111111111111111110011111111111111111111111111110000011111111111111111110000000000000000000011111111111100111111111111111111111111111101111111111110000000000000;
			9'd142: q <= 640'b0111110000000000000000000000000001100011101111110000111111111111111111110100100000000000000111111111110000000000000001111111100000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000001100000000000001111111111111111111111111111111111111111111111111111110000000000000000000000000000000011111111111111111111111111111111111110011111111111111111111111111111111111111111111110011111111111111111111111111110000011111111111111111100000000000000000000001111111111100011111111111111111111111111111111111111100000000000000;
			9'd143: q <= 640'b1111110001000000000000000000000001000011101111100000111110101001011011111100100111001111111111111111111000000000000000111010000000000000000010110000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000011100000000000001111111111111111111111111111111111111111111111111111110100000000000000000000000000000011111111111111111111111111111111111110111111111111111111111111111111111111111111111110011111111111111111111111111110000011111111111111111100000000000000000000001111111111100111111111111111111111111111111111111111100000000000000;
			9'd144: q <= 640'b1111111000000000000000000000000011000011101111000001111110010011111111111100100111111111111111111111000000000000000000000000000000000000001000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000011100000000000001111111111111111111111111111111111111111111111111111111100000000000000000000000000000011100011111111111111111111111111111110111111111111111111111111111111111111111111111110011111111111111111111111111000000011111111111111111100000000000000000000001111111111100111111111111111111111111111111111111111000000000000000;
			9'd145: q <= 640'b0101111000000000000000000000000000000001101111000001111110011111111111111100101011111111111111111110000000000000000000000000010000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000011000000000000001111111111111111111111111111111111111111111111111111111100000000000000000000000000000011000001111111111111111111111111111110111111111111111111111111111111111111111111111110011111111111111111111111111110000011111111111111111100000000000000000000001111111111100111111111111111111111111111101111111111000000000000000;
			9'd146: q <= 640'b0111110000000000000000000000000000000001100111010001111111111111111111111100000011100011110110111110000000000000000000000000010000000000000001011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011000010000000000000001111111111111111111111111111111111111111111111111111111100000000000000000000000000000011000001111111111111111111111111111110111111111111111111111111111111111111111111111110011111111111111111111111111110000011111111111111111100000000000000000000001111111111100111111111111111111111111111101111111110000000000000000;
			9'd147: q <= 640'b1111110000000000000000000000000000000001100111000001111111111111111111111100000111111000111101111010000000000000000000000000001000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000001111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000001111111111111111111111111111110111111111111111111111111111111111111111111111110011111111111111111111111111110000111111111111111111100000000000000000000011111111111100111111111111111111111111111111111111110000000000000000;
			9'd148: q <= 640'b1100000000000000000000000000000000000001100111010001111111111111111111111100000101000000011100001000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000001111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000001111111111111111111111111111110111111111111111111111111111111111111111111111110011111111111111111111111111110000000001011111111111000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000;
			9'd149: q <= 640'b0000000000000000000000000000000000000001110111000000000000011111111111111100111111111111011101011100000000000000000000000000000100000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000011111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000001111111111111111111111111111100011110000000000000000110000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd150: q <= 640'b0000000000000000000000000000000000000001110010000000000000111111111111111100111111111111111111111111000000000000000000000000001110000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000111111111111111111111111111111100111111001111111111111000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd151: q <= 640'b0010000000000000000000000000000000000001110011000000000000111111111111111100111111111111111111111111000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd152: q <= 640'b0011010000000000000000000000000000000011110011000000000000011111111111111100011111111111111111111111100000000000000000000000010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd153: q <= 640'b0011100000000000000000000000000000000011111011000000000000011111111111111100011111111111111111111111100000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd154: q <= 640'b1001000000000000000000000000000000000011011111000000000000001111111111111100111111111111111111111111100000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd155: q <= 640'b0100100000000000000000000000000000000011100011111000000000001111111111111100111111111111111111111111111100000000000000000001000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd156: q <= 640'b0000101000000000000000000000000000000011111000000000000000001111111111111100111111111111111111111111111111000000000000000000100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000111111111111111111111111111111111111110000000000000000000000000000000111111111111111011111111111111111011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd157: q <= 640'b0000000000000000000000000000000000000011110000000000001000000111111111111100111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000000000000000000000000000001011111111111111111111000011111111111111111110000000000000000000000000000111111111111111111110011011011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000;
			9'd158: q <= 640'b1111110000000000000000000000000000000111110111100000001100000111111111111110011111111111111111111111111001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000011111111111111111111111111111111111111111111111110000000000000000000000000000111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd159: q <= 640'b1111100000000000000000000000000000000000111111110000000100000011111111111100011111111111111111111111110001100000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000100000000111111111111111111111111111111111111111111111111110000000000000000000000000000100111111111111111111111111111111111111011000111111111111111111100000000000001000000000000011111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000;
			9'd160: q <= 640'b0110000000000000000000000000000000000000000000000000000001100011111111111110111111111111111111111111001000100000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000001110000111111111111111111111111111111111111111111111111111110000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111100000000001111111111000000000000000000000000000000000000000000000000011111111110000111000000000110000000110000000;
			9'd161: q <= 640'b1111000000000000000000000000000000000000000000000000000001000011111111111110011111111111111111111110000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000001110000111111111111111111111111111111111111111111111111111110000000000000000000000000011111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111011111111111111111111111111000000011111111111111111111111100000000000000011111111111101111111111111111111111111111111111111110000001111000000;
			9'd162: q <= 640'b0001000000000000000000000000000000000000000000000000000010000001111111111110011111111111111111110110010000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000001110000111111111111111111111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111011111111111111111111111111000000111111111111111111111111100000000000000011111111111101111111111111111111111111111111111111110000001111000000;
			9'd163: q <= 640'b1000000000000000000000000000000000000000000000000000000010000001111111111110011111111111111111001010000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000001110000111111111111111111111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111011111111111111111111111111100000011111111111111111111111000000000000000011111111111101111111111111111111111111111111111111110000000111100000;
			9'd164: q <= 640'b1111000000000000000000000000000000000000000000000000000010000000111111111100011111111111111110000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000001100000000000000001111000111111111111111111111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111100000111111111111111111111111110000000000000011111111111101111111111111111111111111111111111111110000000111110000;
			9'd165: q <= 640'b0100000000000000000000000000000000000000000000000000000001000000111111110100011111111111001110000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000001100000000000000001111000111111111111111111111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111100000011111111111111111111111110000000000000011111111111101111111111111111111111111111111111111111000000111110000;
			9'd166: q <= 640'b1111000000000000000000000000000000000000000000000000000000000000001111110010011001101000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000000000000000001100000000000000001111000111111111111111111111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111000000011111111111111111111111111000000000000011111111111111111111111111111111111111111111111111111000000111110000;
			9'd167: q <= 640'b1111001000000000000000000000000000000000000000000000000000000001111110001000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000001100000000000000001111000111111111111111111111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111100000011111111111111111111111111000000000000011111111111101111111111111111111111111111111111111111100000011100000;
			9'd168: q <= 640'b0110000000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000011000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000001100000000000000001111000111111111111111111111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111011111111111111111111111111100000011111111111111111111111111000000000000011111111111101111111111111111111111111111111111111111110000001100000;
			9'd169: q <= 640'b0100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000001010001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000001100000000000000001111010111111111111111111111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000111111111111111111111111111000000000000111111111111101111111111111111111111111111111111111111111000000000000;
			9'd170: q <= 640'b0100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000100000000000000001111000111111111111111111111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111111111111111111111111111000000000001111111111111101111111111111111111111111111111111111111111100000000000;
			9'd171: q <= 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000100000000011000001111111111111111111111111111111111111111111111111111111111110000000000000000000000000111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111110011111111111111111111111111000000011111111111111111111111111000000000111111111111111111111111111111111111111111111111111111111111110000000000;
			9'd172: q <= 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000011111111100000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000100000000000000001111110111111111111111111111111111111111111111111111111111110000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111000000011111111111111111111111111000000001111111111111111101111111111111111111111111111111111111111111110000000000;
			9'd173: q <= 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000011100011111111110000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000001111000111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111110000000011111111111111111111111111000000011111111111111111101111111111111111111111111111111111111111111111000000000;
			9'd174: q <= 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000011100011011111111000000000001000001111111110111111111111111111111111111111111110000000000000000000000000000000000000000000000000111100000000000000000000000000100000000000000001111010111111111111111111111111111111111111111111111111111111000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111110000000011111111111111111111111111100000011111111111111111101111111111111111111111111111111111111111111111000000000;
			9'd175: q <= 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111100000000000000000001110000111111111100000000000000000000000000000100000000000000000001000000000000000000000000000000000000000000000010111111100111111100000000000000000111111111101111111100000001111010111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111110011111111111111111111110010000000011111111111111111111111111100000111111111111111111111111111111111111111111111111111111111111111111110000000;
			9'd176: q <= 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000111000111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000010001100000000000000001111000111111111111111111111111111111111111111111111111111111100000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111000100000000011111111111111111111111111000000011111111111111111111111111111111111111111111111111111111111111111110000000;
			9'd177: q <= 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100001111000000000000000000111000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111000000000000000000000000001100000000000000001111000111111111111111111111111111111111111111111111111111111100000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111100000000011111111111111111111111111000000011111111111111111111111111111111111111111111111111111111111111111110000000;
			9'd178: q <= 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000111000000000000000000011000001111111111000000000011000011100000001110000000000000000000000000000000000000000000000000000000000000000000000000000011010000000000000000000000000000100000000000000001111000111111111111111111111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111101110011111111000000000000011111111111111111111110111000000111111111111111111111111111111111111111111111111111111111111111111110000000;
			9'd179: q <= 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000011000000000000000000011100001111111111100000000000000000000000001111111111111111100000010000000000000000000000000000000000000000000000000000000011000000000000000000000000000000100000000000000001111000111111111111111111111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011110011000101100010000000000000001111111111111111111110111100000111111111111111111101111111111111111111111111111111111111111111111110000000;
			9'd180: q <= 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000010000000000000000000011110000111111111110000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000001111000111111111111111111111111111111111111111111111111111111110000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111010000111100101100000000000001111111111111111111110111100000111111111111111111111111111111111111111111111111111111111111111111100000000;
			9'd181: q <= 640'b0000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000001111111111111100011000000000000000000001110000111111111110000000000000000000000000011000100001000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000001111000111000111111111111111111111111111111111111111111111111111000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111110011111111111110000000000001111111111111111111110111000000111111111111111111111111111111111111111111111111111111111111111111100000000;
			9'd182: q <= 640'b0000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000001111111111000010111000000000000000000001110000111111111111000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000001111111111111111111111111111101111111111111111111111111000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111110111111111100000000000000011111111111111111111110111111000111111111111111111101111111111111111111111111111111111111111111111000000000;
			9'd183: q <= 640'b0000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000010000000000001111110000001111000000000000000000000111000111111111111000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000011010000000000000111111111111111111111111111111001111111111111111111111111000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011101111000111110000011000000000011111111111111111111110111100000111111111111111111101111111111111111111111111111011111111111111111000000000;
			9'd184: q <= 640'b0000000000000000000000000000000000000011000000000000000000000000000000000000000000001000001111010000000000000000001111110000001111100000000000000000000111100011111111111100000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000011111111111111111111111110001111111111111111111111111111000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111110000000000000000001111111111111111111111111100000011111111111111111101111111111111111111111111111111111111111111110000000000;
			9'd185: q <= 640'b0000000000000000000000000000000000000010000000010000000000000000000000000000000000111111111010000000000000000011111111111100000111100000000000000000000011100011111111111100000000000000000000000000011111111110000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000111110111111111111111111111100110111111111111111111111100000000000000000000011111111111111111111111111111111111111111100111111111111111111111111111111111111111111111110011111100000001100000000000000000000111111111111111111101111000000011111111111111111101111111111111111111100000000000000000000000000000000000;
			9'd186: q <= 640'b0000000000000000000000000000000000000010000000010000000000000000000000000000001111111111100010000000000000100111111111111101111111100000000000000000000011100001111111111110000000000000000000111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000001111111111111111111111111111101111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000011111110000000000000000000000000111111111111111100111111000000001111111111111111111111111111111111110000000000000000000000000000000000000;
			9'd187: q <= 640'b0000000000000000000000000000000000000000000000000000000000000000000001111110000000100000110110000000000000001111111011111111111111100000000000000000000011110010111111111111000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000011111111111111111111011111111101111111111111111111111000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111100111110011111111111111111110001111111100000000000000000000000011111111000000000011000000000001111111111111001111111111100000000000000000000000000000000000000000000;
			9'd188: q <= 640'b0000000000000000000000000000000000000000000000000000000000000001111111000000000000111100010000000110000001011111110011111111111111100000000000000000000001110000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000111111111111111111111111111111111111111111111111111111000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111110000111111111000000000000000000000000000000000000000000000000000000000000000000000011110100000000000000000000000000000000000000000000;
			9'd189: q <= 640'b0000000000000000000000000000000000000000000000000000000011111110000000000000000011111111010000110110010110111110000011111111111111100000000000000000000001110000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000111111111111111111111111111111111111111111111111111000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100101110000011111111110000000000011111111110000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000;
			9'd190: q <= 640'b0000000000000000000000000000000000000000000000000000001111000000000000000001011111111111111111111111111111111100000011111111111111100000000000000000000000110000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001111111111111111111111111111111111111111111111111111000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011011111111000001111111100000000011111000000000000000000000000000000000111100001111111110000000000000000000000000000000000000000000000;
			9'd191: q <= 640'b0000000000000000000000000000000000000000000000100000000000000000000000001111001111111111111101111111111111111100000111100101111111100000000000000000000000111000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000011111000000000000001111111111111111111111111111111111111111111111111111000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111101111000000000111111111100000001000000000000000000000000000000111110001111111111111110000000000000000000000000000000000000000;
			9'd192: q <= 640'b0000000000000000000000000000000000000000000000000000000000000000010111001111001111111111111111111111111111111000001111100101111111000000000000000000000000111000000111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000001111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111000011011110000000011111111111100000000000000000000000000000000001111001111111111111100000000000000000000000000000000000000000;
			9'd193: q <= 640'b0000000000000000000000000000000001000000000001110000011111111111111111111111001111111111111111111111111111110000001111000101111010000000000000000000000000011000000111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111000000000000000000001101111100111111111111111111111111111111111111111111100000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000100000000011111111111100000000000000000000000000000000000101111010111111000000000000000000000000000000000000000;
			9'd194: q <= 640'b0000000000000000000000000000000000100000000000000000011111111111111111111111111111111111111111111111111111110000000111000001111000000000000000000000000000011000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000001111010111111111011111111111111111111111111111111111100000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111110000111111111111100000000000000000000000000000100000000111011100000000000000000000000000000000000000;
			9'd195: q <= 640'b0000000000000000000111111000000000100100000000110000011111111111111111111111011111111111111111111111111111100000000010000000110000000000000000000000000000001100000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000001111111110001111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110001111111111111000000000001000100111101100001111110000000000000000000000000000010111111100000000000000000000000000000000000000000000;
			9'd196: q <= 640'b0000000000111111110000000000000001000000000000110000011111111111111111111111111111111111111111111111111111100000000000000000010000000000000000000000000000000110000001111111111100000000000001000000001100010000000110111100000000000000000000000000000000000000000000000000000000000000000000000001111111000111111111111000000000000000001111111111111111111111111111111111111111111111111111000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001000000010000000000000000000110010111111111100000000000000000000000011111111100000000011111110000000000000000000000000000000000000000000;
			9'd197: q <= 640'b0000111111100000000000000000000000000000000000110000001111111111111111111111111111111111111111111111111111000000000000000000000000000001100000000000000000000110000000011111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000111001111111110110000000000001111111111111111111111111111111111011111111111111111110000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111100000000000000000000010000000110011111111110000000000000000000000000001111111111111111100000000000000100000000000000000000000000000000000;
			9'd198: q <= 640'b1111111111111111111111111000000000000000000000000000000111111111111111111111111111111111111111111111111110001100000000000000000000000011000000000000000000000011000000001111110000000001111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000010000001111111111111111111111111111111111111111111111110000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110000001000000000000000111111111010000000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000;
			9'd199: q <= 640'b1000000000000000000111111111111100000000000001110110000011111111111111111111111111111111111111111111111111011110000000000000000000000011000000000000000000000111000000001111111000000000000000000000000000000000000000000000000001111000011110000111111100111000000000000000000000000001111000000000000000000000100000000000000001100000000111111111111111111111000001111111111111111111111110000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011110001100001000000000000000000111000000000000000000000000000000000000000010000000000000111111111111110000000000000000000000000000000000;
			9'd200: q <= 640'b0101101010000000000000000000000000000000000000100000000001111111111111111111111111111111111111111111111111111100000000000000000000000001010000000000000000001111000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100000001100000000000000000000000000110000000010110000000000001111111111111101100000001111111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100101111100100001000000000000000000000000000000000000000000000000000000000000000000000010000000000001111111111111111100000000000000000000000;
			9'd201: q <= 640'b1100000000000000000000000000000000000000000000000000000001100111111111111111111111111111111111111111111111111100000000000000000000000001111110000000000001111111100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000111110000000000000001111111111111110000011111111111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001111111110010000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110000000000000000000;
			9'd202: q <= 640'b1101100001000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000001111111111111111111111111111111111111111111111111100000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111001001011111111010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd203: q <= 640'b1111111100000000000000000000000000000000000000000000000000000011111111111111101111111111111111111111111110000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000111111000011111111111111111111111111101111111111000000000000000000000000000101111111111111111111111111111111111111111111111111111111111111111111111111111111000001111111000011111110110011000000110000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd204: q <= 640'b1101111011111111001111001100000000000000000000000000000000111111111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000001000000000000000000111111100000000000000000000000000000000011111111111111111111111111111111111111001000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111110110011111111110000000110000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd205: q <= 640'b1111111111111111111111000100000000000000000000000000011001111111111111111111111111111111111111111111111100000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000001111000010111100000000000000111111000000000000100000000000000000001111111111111111111111111111111111111111111111000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111010010111111111101100001101000000000000000000001000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000;
			9'd206: q <= 640'b1111111111111111111111110000000000000000000000000000000000011111111111111111111111111111111111111111111100000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000111111000000000000111110000011100000000000000000000000001111111111111000001111111110000011111111111111111000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000111010001100000000111110011111111000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000;
			9'd207: q <= 640'b1111111111111111110111001000000000000000000000000000000001111111111111111111111111111111111111111111111100000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000001110000111111100000001111100000000000000000000100000000000000000111111110000001111100000001111111111111111101010000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111110001100000101101011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd208: q <= 640'b1111111111111111111111111110000000000000000000000000000111111111111111111111111111111111111111111111111100000000000000000000000000000000000001111111111111111111110000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000001110000001111000011111000000000000011111111111110000000000000001111110000000000000111111111111111111000111111110000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100111101111111111111110000000000001111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000;
			9'd209: q <= 640'b1111111111111111111111111111000000000000000000000000000111111111111111111111111111111111111111111111111110000000000000000000000000000000000011111111111111111111100000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000000100000111111111110000000000111011111111101000000000000000000000000000111111111111111111000000111111111111111110000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111100011111110111111111111000000000000001001110000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000;
			9'd210: q <= 640'b1111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111000000000000000000000000000000000011111111111111111111100000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000110000111111100000000000000000000000000000000000000000000000011111111111111110000010011111111111111111000000010000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111000000001100111111100000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000;
			9'd211: q <= 640'b1111111111111111111111111111111000000000000000000000001111111111111111111111111111111111111111111111111111100000000000000000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000001000000000000000000111111111110000000000001111111111111111111111111111111110000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111110100000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000;
			9'd212: q <= 640'b1111111111111111111111111111111111111111000000000000011111111111111111111111111111111111111111111111111111100000000000000000000000000001000111111111111111111111100000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111100000000000000000000000000000111111111100000000000000010000111111111110001111111111100011111111110000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000100000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000;
			9'd213: q <= 640'b1111111111111111111111111111111111111111111111111000011111111111111111111111111111111111111111111111111111110000000000000000000000000010000111111111111111111111100000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000001111110000111111100000000000000011111111111111000000000000000000000000000001001111010101111111111111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111110000001100100000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000;
			9'd214: q <= 640'b0001111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111100000000000000000000000000000111111111111111111111000000000000100000000000000000000000000000000000000111110000000000000000000000000000000000000000000011111110000000111111100000111111111111000100000000000000000000000000000000000000111111111111111111111111111001111111111000000000000000000000001111111111111111111111111111110111111111111111101111111111111111111100000101001000001110001111000001111110111000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000;
			9'd215: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000111001111111111111111111111000000000000000000000000000000000000000000000001110001111111100000000000000000000000000000000000011111000000000111111111111110000000000000000000001100000000000000000000000000100001111101111111111111111111111111111111101000000000000000000000000111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000;
			9'd216: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111111111111111111111111110000000000000000000000000000000010011111111100000100000000000000000000000000000000000000000001111111000001111111111111111000000000000000000000000100000000000000000000000000000000011111111111111111111111111111111111111110000000000000000000000000111111111111111111111111111111111111111111111111111111111111111110100111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000;
			9'd217: q <= 640'b0001100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111110000000000011111000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000001111111111000000000000011110100000000000000000000000000000000011111111111111101111111111111111111100111010110000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111000111111000000010000000111111101111111111101100000000000100000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000;
			9'd218: q <= 640'b1111111110000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010000000000000001000000111111111111111111111110000000000011100000000000000000000000000000000000000000000000000000011111111111100000111111000000000000000000000001111111100000000000000111111111111111000000000000000000000000011101111111111111111111111111111111111111101101111111000000000000000100111111111111111111111000011111111111111001111111111111111111111110011111110011100000011111100000000000000000000000000000001100000000000001111110000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000;
			9'd219: q <= 640'b0011111111000000111011010001111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000001111111111111111111111111111110000000001111110000000000000000000000000000000011111111111111111110000000000000000011110000000000000000000011111111111110000000000000000000000001001100000000000000000000001111111111111111111111111111110111111111011111100000000000000000000000000000011111111111111111100011111111111111110011111111111111111111100011111110000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111101000001111100000000000000000000000000000000000;
			9'd220: q <= 640'b0011111111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111100000000100000000001111111111111111111111111111110000000001111110000100000111111111111111111111000000000000000000000000000000001111100000000000000000000000011111111101000000000000000000000000000100000000000000000000000000011111111111111111111111111111111111111110000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111110001111000000000000000000000000001000000000000000010000000000000001000000000000000000000000000000000000001000001001111111111111111100111000000000000000000000000000;
			9'd221: q <= 640'b0111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111110000000000011000000000111111111111111111111111111110000000011111111111111111111110110000000000000000000000000000000000000000011111000000100000000000000000000011110000001111100000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111010000000000000000000000000000111111111111111111111111111111111111111111110111111111111110110101000001111000000000000000011110010000000000000000110111000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000;
			9'd222: q <= 640'b1111111111111111110000000000000000101111111111111111111111111111111111111111111111111111111111111111111111100000000000011111000000000001111111111111111111111110000000011111110000000000000000000000000000000000000000000000000000000111110000000000100000000000000000000011100001111111100000000000000000000000000000000000000000000000000001111111111111111111111011110001111111011111111110000000000000000000000000001111111111111001111011111110111111111110100110110111111010111110000000111000000000000000001000000000000000000000000110100000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000;
			9'd223: q <= 640'b1111111111111111111000000000000000010111111111111111111111111111111111111111111111111111111111111111111111000000000000011111100000011111111111111111111111111111000000111111110000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000000110011111111111111101010000100000111010000000111000000000001100000000000001111111111111111111111111111111100000010000000000000011111111010000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000;
			9'd224: q <= 640'b1111111111111111111100000000000000000111111111111111111111111111111111111111111111111111111111111111111111000000000000011111110001111111111111111111111111111111110000011111100000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000011111111011111100000000000000000000000000000000000000000000000000000010111111111000100000000000011111100000010010000000000000111111111110110000000001111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000;
			9'd225: q <= 640'b1111111011111111000000000000000000000000001101101011111111111111111111111111111111111111111111111111111110000000000000011111100011111111111111111111111111111111111100011111100000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000000000001111100000110010000000000000010111011111111100000000000000000000000000000000000000000001001110000000011011011111111111111111111111111111111111100000000110000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000;
			9'd226: q <= 640'b1111111111111111111111110000000000000000000000001000010001110111111111111111111111111111111111111111111111000000000000011111100011111111111111111111111111111111111110100111100000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000011111110000000000000000000000000000011100000000000000000000000000010000000000000000000000000000001111111111101110000000000000000000000000000000000000101111111100000110111001000000000111111111111100111111111111111111111111111111001000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000100000000000000000000;
			9'd227: q <= 640'b1111111111111111111111111111110000000000000000000000000000000011111111111111111111111111111111111111111111100000000000011111100000011111111111111111111111111111111111111111000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000001100000001000000000000000011111100011111111100000000000000100000000000000000010100001111101110000011111111100000011110000110111010000010000000000011111111000111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000001110000000000000000000;
			9'd228: q <= 640'b1111111111111111111111111111111010000000000000000000000000000001111111111111111000011111111111111111111100000000000000111111000001111111111111111111111111111111111111111100000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000110010011000000000001111111111111111111111111110000000000000000000000000001111110000001111110000001111011111000000110110000111101111111111110100000000000000000000000000000000111111111111111111111111111111011111000000000000000000000000000000000000000000000111111000000000000000000000000011100000000000000000000;
			9'd229: q <= 640'b1111111111111111111111111111000000000000000000000000000000000000011110111111111000001111111111111111111100000110000001111111100011111111111111111111111111111111111111111110000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011100001111111111111111111111111111111111110000000000000000000000000011111100001111111000000001011111100001101111000000000000111111111110000000000000000010000000000000111110000000000000000000000000000111111111111100000000000000000000000000000000000011111100000000000000000000001111111110000111000000000000;
			9'd230: q <= 640'b1111111111111111111111111111111111111111100000000000000000000000000010111111101000001111111111111111001111111000000001111111100011000011111111111111111111111111111111111110000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111111111111111111111111111111111111110000000000000000000000000111101001111111100000000111111111100011111001000000000000110011000010000000000000000000000000000100111111111100000000000000000000000000000000000000000000000000000000000000111111110111111000000000000000000000111111111111000111110000000000;
			9'd231: q <= 640'b1111111111111111111111111111111111100111111111110000000000000000000001001111001000000111111111111000000000000000000001111111000000000001111111111111111111111111111111111110000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000111111111111111101011111111111111110000000000000000000000000111111111111111001100001111111111100000100000000000000001100000001000000000000000000000000001000010000111111000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000111100111001111111110000000000;
			9'd232: q <= 640'b1111111111111111111111111111101000000000001111111110000000000000000000000000000000000011111111110000000000000000000001111110000011111101111111111111111111111111111111111111000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000011111111111100001111111111111010000000000000000000000000000111101111111110111111011111111110010001101000000000000000010000000000000000000000000000000000000000001111111000001100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000111000000111111111110000000000;
			9'd233: q <= 640'b1111111111111111111111111110111111110000111111111111111000000000000000000000000000000001111111111000000000000000000001111100000011111111111111111111111111111111111111111111000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000111111111111111111111111111111100110000000000000000000000000000111111111111111111111111111101110101011111111111111000000000000000000000000000000000000000000000111111111001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000111111111111000000000;
			9'd234: q <= 640'b1111111111111111111111111111111111100011111111111111111111010000000000000000000000000000111111111000001110000000000011111100000011111111111111111111111111111111111111111111001100001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111110111110000000000000000000000000111100111111011111111111110000110111111111111111111001000110100000000000000000000000000010110000100011110000011000000100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111101111111111110000000000;
			9'd235: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111011100000000000000000000011111111000001110000000000011111100000001100011111111111111111111111111111111111111100011111111000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111011111111111111111111111111111111000000000000000000000000000000001111111111111111111110000111111111111111111111100011111111110000000000000000000001110000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000111000000000000000000;
			9'd236: q <= 640'b1111111111111111111111111111111111111111111110111111111111111111111111110000000000000000001111111000000000010000000011111100000011111111111111111111111111111111111111111111111111110000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111001111111111111110111000000000000000000000000000000000111111111111111010011000011111111111111111111100111111100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000;
			9'd237: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000011111000000000000000000001111000000011111111111111111111111111111111111111111111111100000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010000000000000000011110001010000000110011000011000000110011000001100000000000000000000000000000000110111110000111001100000001111111111111111111111000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000;
			9'd238: q <= 640'b1111111111111111111111111111111111101111111111111111111111111111111111111111111000000000000001111000001110000000000011111000000011100001111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000111111110011100000011111111111111010011111110000000000000000000000000000000000000001110000000011111110000010000110011111111111111111110000000000000000000000011111010000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000;
			9'd239: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000011010000111000000000011111000100010000000111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000001000011111111111111111111111111111110100000000000000000000000000000000000000000000001111000000000111110010011111111000000011101000001000000000000111011001101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000;
			9'd240: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000011100000011110000000011111000000000000001111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000011111111111111111000111111111111111110011100000000000000000000000000000000000000000000000000001000110000000101111111000000000000101110000000000011110101111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000;
			9'd241: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111100000000000000000011111000100001101001111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111101111111111111111100100000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000011111111101111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000;
			9'd242: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011100000000000111110000000001000001111111111111111111111111111111111111111101100000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000001001111111101111111110000111111111111111100011100000000000000000000000000000000011000000000000010000000000000000000000000000000001110000000001111110000000001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000;
			9'd243: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111000000001111110000000001100000111111111111111111111111111111111111111111111110000000000000000000000000100111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000110000011111111111111100011111111111111100111110000000000000000000000000000000001100000000101001111110100000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000;
			9'd244: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011000000011111110000000000000000111111111111111111111111111111111111111111110000000000000000000000000000000000000000000001111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100111111111111111001011111111111111111000011110000000000000000000000000000001110000000000000011111011000000001111110000100000011000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd245: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000011111110000000000000000111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000111000000011111100011111111111111100001111111000000000000000000000000000000000000000111111111011111000100111111110000000000000000000000011010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd246: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111110000000000000000111111111111111111111111111111111111111111111001000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000100000000000000000000001000000000000000000000000000011111111111011111111110000000000000000000000000000000000000000111111111111110000101111011000000000000000000000000000000000000000000001111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd247: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111000000111111100000000000000000111111111111111111111111111111111111111111111100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111000000000000000000000000000000000100001101111000000000100000000000000000010000000110111101110001000000000000000000000000000000000000011111111111100011111110001101001000000000000000000000001111000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd248: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111000000111111110000000000000000111111111111111111111111111111111111111111111110101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000001111111111000000111111100000001111111100000000000000000000110000000000000000000000000000111111001111111111111100010001111111110100000000000000000000000011111000000000111001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd249: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000111111110000000000000000001111111111111111111111111111111111111111111111111100000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111110000000000000001111111111111111111111111111000000000000000000000000000000000000000000000111100001111111111111111111111111111100100000000001000000000001111100000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd250: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000111111110000000000000000011111111111111111111111111111111111111111111111000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111110000000000000011111111111111111111110111100111011000000000000000000000000000000000011111111111111111111001111111110100000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd251: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111111110000000000000000011111111111111111111111111111111111111111111000000000000110000000000001000011000010000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000001111111111111111111111111111110000000001111110111111111111110000000000000000000000000000000000000000000000000111111111111111100000000010011000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd252: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000010000000111111111000000000000000011111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000110011111111110000000000001111111111111111111111111111000000001111111111100000000000000000000000001000111100000000000000000000000001011000000000000111000000010000000000011010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd253: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000001111111111000000000000000001111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000111111111110111111110000000000001111111111111111111111111111100000000000000000000000000000000101111111111111111110100000000000000000000000000000000000000000000000000110000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd254: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000001111111111000000000000000001111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000001111000000000011111110111111111111111100000000000111111111111111111111100000000000000000000001111111111111111111111111000111100000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd255: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000110000000111111111111000000000000000001111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000001100000000000000001000001111111111111111111111111111111111101000000000001111111111111111111000000000000000000001101111011111110011111000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd256: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000111111111111100000000000000001111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000001111000000000000000000110111111111111111111111111111111111111111111111111111101000000000000000000001111111111111111111111111000000000001100001000111100000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd257: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111111111111100000000000000001111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000010111111111111111111011111111111111111111111111111111111111111100000000000000000000000001111111111111111111111111111000000000000000000000001101100011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd258: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111111111111100000000000000000111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001111000000000111111111111111111111111111111111111111111111011111111111110000000000000000000000000000000000000000011111111111111111111111111111100000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd259: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000001111111111111110000000000000000111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000111100000000111111111111111111111111111111111111111111111111111111111111110000000000000000000000000001111111111111000000000000000001111111111111111111111111111000000000000000000000000100000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd260: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111110000000000000000011111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000100111001000000000000111101110111111111111111111111111111111111101111111111111111111100000000000000000000000000111111111010000001111111111100000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd261: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111110000000000000000011111111111111111111111111111111111111111100000001100011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000001110000111100000000000111111111111111111111111111111111111111111111111000000000000000000000000000011100100000000011111111110000011111111000000000000000000001111111111111111111111111000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd262: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111000000000000000011111111111111111111111111111111111111111100000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000111110000000000000000000000011111111110001110111111111111100111111000000000000000000000000000000010000000011111111111000001111111111100000000011100000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd263: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000001111111111111111000000000000000001111111111111111111111111111111111111111111000000000000000000000000000000000001111111111111111100000000000000000000000000000000000000000000000000000000000000000001111100000111100000000000000000000000011111111110011111111111111111111111111100000000000000000000000000000000011111111111111111100000010001111110000000000000000000000111111110000000000000000000011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd264: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111000000000000000001111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000011000001100000000000000000000000000000111111111111111111111111111111111110000000000000000000000000000000000111111111111111111100000000001111000000000000000000000000000000000000000000100000000000000000000000011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd265: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111100000000000000000111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000011000110000000000000000000111111111110111111111101111111111111010111111111000000000000000000000000000000000001111111111111111100000000001111110000000000000000000000000000000000000000000000000000000010000100000000000000000000011111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd266: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111100000000000000000111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000011001010000000000000000000001111111111111111111111101111111111101011111111111010000000000000000000000000000000011111111111111111000000000000000111111000000000000000000000000000000000100000001000011000000000000000000000000000000000000000000000001111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd267: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000011111111111111111110000000000000000111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000001111110000000000000000000001001100111111111111111111111111111111111111111111110000000000000000000000000000001111111111111111100001000000000000111110000000000000001110000000000011001000000000001111000001000000000000000000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000000000000;
			9'd268: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000011111111111111111110000000000000000111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000001100000011110111111111110111111111000001111111111110010111100000000000000000000000000011111111111111111100100100000000111100000000000000000000010000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111110000000000000000000000000000000000000000000000;
			9'd269: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000011111111111111111110000000000000000111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000001111111111111110011011111111110001111111111111111111111100000000000000000000000000011011111111111100000001000000010111000000000000000000001111011100000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000;
			9'd270: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111111111111111111110000000000000000111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000111101111110001111111111111111111111111000000000000000000000000000000000111111111000011110000011111000000000000000000001011111111111101111110000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000;
			9'd271: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111000000000000000011111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011111111111111111111100000000000100000111111111111111111111111011000000000000000000000000000000000000111000001110000000111111000000000000000000000000000110111000010000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000;
			9'd272: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111000000000000000011111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000011111111111111111111110000000000001111111111111111111000000000000000000000000000000000001100000000000000001101111000000000011110100000000011110100000000000100000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111;
			9'd273: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111111111111111111111000000000000000011111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100001111111000000000000000001111111111111111111111111100000111111111111000000000000000000000000000000000000000010110000100000100111000000000000110000000000111110111000000011000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd274: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000001111111111111111111111100000000000000011111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000001111111111111111111111110000000000000000000000000000000000000000000000000111101110011111111110000000001000000001100000000100000001110000001000000000000001100000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd275: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000001111111111111111111111100000000000000011111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000111111111111111111111110000000000000000000000000000000000111100111111111111101000000000000000000000111100000110000000111100000000000000000000111110000000000000110001100000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd276: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000001111111111111111111111100000100000000011111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011111110011000001111111111111100000000001111111111111111110000000000000000000000011111111111111111100010000000000000000000111110000001000000011111000000000000000000001111110000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd277: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111100001100000000001111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000010111110000111111111011111110000000000000000000011111111111110000000000000000011111111010000000000000011000000001111111111110000001111110000000000000000001101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd278: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000011111100000011010101101000011111111111000000000000000000010111111111111111110000000000000110001000000000000000111111111110000000111100000000000000000000011011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd279: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001100000000001111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001111100000000000110000011000000110000000011111111100000000000000000000000000000001111111111111111111111000000000000101111100111110100000000001110000000000000000000000111110011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd280: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000011111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110000000001111100001111001000001100001101110100000000111111111110000000000000000000000000000000000000000111111111111111111111000000000000001100111111000001110000000000000000000111111000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd281: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000111010000111111110000001100001111110000000111111111111010000000000000000000000000000001111101100110000000000011111111111111111111110000000000000001111110000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd282: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000011111111100001111111001111100000011111111110101100000000000000000000000000000001110000011111111110000000000000001111111111111111111111000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd283: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000001110111011100011111001111111111111111111111111111110000000000000000000000000000000000001111001111100000111111111110000000000011111111111111111111111000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd284: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000011011111001000001111111111111111111111111111111111000000000000000000000000000000000000011000000000110010000011111111111110000000000000000011111111111111111111110000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd285: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000111111001000000111011111111111111111111111111111110000000000000000000000000000000000000000000000100000100000011111110000000011110110100000000000000000011111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd286: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000001111111111111111111111111111111111000000000000000000000000000000000000000000000000001000100011111111100000000011111111000000001111000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd287: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111111111000111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000011111101111111111111111111111111111100000000000000000000000000000000000000000000000000100101111111111110000000000011111111100011100000000000001111111110000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd288: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000001111111101111111110101111111110000000000000000000000000000000000000000000000011110001111111111110000000010111111110000001100000000000001110000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd289: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111111111100000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000011111111111111111101111111111111111110000000000000000000000000000000000000000010011111111111111111110110111111111000011000000000000000100000000000000000000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd290: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111111111100000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001101111111111111111110111111111111111111100000000000000000000000000000000000000001100011111111111111111101111111110001111110000000000000000000000000000000000000000000000000000011100000000000000000011111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd291: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000010000000000111111111111111111111111111111111111111111000000000000000000000000000000000000000011000000111111111111111111111111000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd292: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000011111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000111111111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111110000000000000000000000000000000000000000001111111111111111111110111111111111100111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000001111000000000000000000000000000000000000000000000000000000000000;
			9'd293: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000011111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111010000000000000000000000000000000000000000001111111111111111111110000000001111111100000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001111111111111111100000000000000000000000000000000000000000000000;
			9'd294: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000011111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000111111111110111111111111111111111111111100111000000000000000000000000000000000000000011111111001100111110111100100000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111110000000000000000000000000000000000;
			9'd295: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000110000111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111000000000000000011000000000000000011111111111111111111111111111111000000011101111000000000000000000000000000000000000000011111111100000111110111100010111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111100000000000000000000000;
			9'd296: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000001110000111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000001111111111111111111111111111111100000000001111100000000000000000000000000000000000000000111111111101000111110111111001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000000000;
			9'd297: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000011110000111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000111111111111111111111111111111111000000010001111010000000000000000000000000000000000000000110000000000011111100111111110000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100;
			9'd298: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000011111001111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111100000000111111111111111111111110000000100000001000000000000000000000000000000000000000000110000000000001111000111111110000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111;
			9'd299: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111011111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111100000000111111111110111000010000111111000000000000000000000000000000000000000100001100000000000111111111111100000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd300: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111110000000010111111101011111111110000000000000000000000000000000000000000001100000000111111111111000100000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd301: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111101000000000001111111111111111111100000000001111111111111000000000000000000000000000000000000000101000000001111111111111101100000000011111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd302: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000111111111111111111110000000101111100000000000000000000000000000000000011111000000011001111111110101111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd303: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000001111111111111111111111000000000000000000000000000000000000111111111000001111111111111110101011100011111111100000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd304: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000001100000000000000000000000001111111111000000000111111111111111111000000000000000000000000000000111111100000001111111111111110101111101111000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd305: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000001111111111100111100000000001111111111111111111100000000000000000001111110000000011111111001111001100111001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd306: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000011111111110000100011111111111100000000001111111111111111100000000000011100110000111110111111111111111001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd307: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000001111110000000000111111111111111111000000000000000011111111111111111100000000001111111111100111111111001000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd308: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000011111000000000011111111111111111110011100000000000000000000111111111111111111100000000001111011111100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd309: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000001111111110010001001000111100000000000000000000000000011111111111111111111110000010000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd310: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100111111111000111100100011111111000000000000000000000000100000000011111111111111111111111000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd311: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000011111111100111111101111111111000000000000000000000000000011111111000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd312: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000011111111111111000000000000000000000000000110111111111111000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd313: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011111011111111111110000000000000000001111111111110000000000000000000000000000111111111111100000000000100000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd314: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111111111111111111111000000000000000000000000000000000000000000000000000111111111000000000000000000011111000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd315: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000011110000000000000000000000000000000000000111111111110000000000000110000111110000011001110000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd316: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000111111000000001111111111111101000000000000000000000000011111111111100000000000000100011111000000000001000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd317: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000111100000000111111111111111111101000000000000000000000000001111111011111000000000000111100000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd318: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000110000000111111111111111110101111000000000000000000000000000000000011111110000000001110000000000000000000000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd319: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000011010001111111111111111110011110000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd320: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000001011111111111111111111111111011110000000000000000000000001000011000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd321: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001111000000000000000000000000111111111111111111111111111111000000000000000000000000100101111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd322: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000001111111111111111111111111111111111000000000000000000000011100000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd323: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100100000000000000000011111111100110011111111111110001000011000000000000000000000000000000000000000100000000110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd324: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001110001100001111111111111111100110001100000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000;
			9'd325: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000010011111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000;
			9'd326: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000011101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000;
			9'd327: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110110111011100000000000000000000000000000000000000000000000000010000100000000111101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000;
			9'd328: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100111111111111101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111110111110011111000111100000000000000000000000000000000000000000010000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000;
			9'd329: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110011111100011000100101100000000000000000000000000000000000001111100000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000;
			9'd330: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111110001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000111111111110111000000000000000000000000000000000000000000000000000000000111111000000111000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000;
			9'd331: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111111110011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000001111111100001101001100000000010000000000000000000000000000000000000000001111110000001101100000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000;
			9'd332: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111100000111111111100011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000001111111000000000000000111100111111000011001111111000000000000000000000000000000000011111111110110111000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111;
			9'd333: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111000000111111111011111111111100111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000011110010110100000000011111111111100000000111111111111000000000000000000000000000000111111111111100100000000001100101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd334: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111100000001111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000001111100111111111010011111111110000000000000000000000000000000011111111111100111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd335: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111000000111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110111110011111111111111111111111110000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd336: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100000111110000101111111100111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000111111111111110111111111111100000000000000011100000000111111111111000010000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd337: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011100001101111000000000111111111111111011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001001000000000000000000000000000000000111111100011111111111000000000000001100000000011111111111110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd338: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000011110011101100000000011111111111111111011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000001100000000000000000000001111111111111100000000000100000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd339: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000011111111001100000000111111111111111110001111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000001110000001111100000000000000000001100111110000000001011000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd340: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000011111111011000011111111110100111111100011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000001110000111000001111100000000000000000000000001111111100000000000010111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd341: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000001111111000001111111111100000000001000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000001111111111000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd342: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000001111111000011111110000000000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000000000111001100001111111111111111111100000000000000000000000000000000000000000000001000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd343: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000001111110001111111100000000000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001010000000000000000111111110001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd344: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000001111110001111111111010000011000110001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000011111111111111111111111111111011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd345: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000001111110000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000011111111011111111111111111111011100101100001100011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd346: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000111110001111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000001111111110111111111111111111111111000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd347: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000001100001111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000011110111110101111111101111100000000000000000011111101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd348: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000011111111111111111111111111111111111111111011100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000110000001100111111111100000000101101111111111010011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd349: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111111111111111111111111111111111111111100000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110000010000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd350: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000001011111111111100000010000000011111000100000000010000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd351: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000111111111111111111111111111111111111111110101111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100111111111111000000001000000011011111100000000000000111110000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd352: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000100000000000000001110101111111111100010100000100000000010011000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd353: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000011111111111000000000001000000000000000000000110001111100000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd354: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000001111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000000100000000000100001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd355: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010110010011110000000000000000000000000000100100011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd356: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000100000000000000000000000001100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd357: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000100000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd358: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000000000000011111111111110111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd359: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000011111111111111111111111111111111111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd360: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000011111111111111111111111111111111111111111011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100000000000000000000000000000001111100111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd361: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000111111111111111111111111111111111111111111111000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000111111111111000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd362: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000111111111111111111111111111111111111111101110001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000011111111111110000000001110000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd363: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000110000000111111111111111111111111111111111111111000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000111110000000011111111111100000000011110000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd364: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111100000000111111111111111111111111111111111111111110111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001110000000001111111111100000000000111000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd365: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001111000000001111111111111111111111111111111111111110111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000010000000000011111111100000000000001110000000000000000110111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd366: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111000000001111111111111111111111111111111111111111111111001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000111111111000000000000110000000000000000001110111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd367: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000100000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd368: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000011111111110111111111111111111111111111111111011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101110100000000000110000000000000000001111011111100001000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd369: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010000001000000011111111101111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000001100000000000011000111111111111100000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd370: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000001111000000111111111111111111111111111111111111111111110000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001000000000000100000000000000001111111111110000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd371: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111000000011111111111111111111111111111111111111111000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001111111111000000000001111000111111111111100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd372: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000110000000011111111111111111111111111111111111111100000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111000000000011111001111111111111000010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd373: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001110000000111111111111111111111111111111111111110000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000001111100011111111111110010000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd374: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001000000000111111111111111111111111111111111111110000000110000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111101111111111110000000011111000011111111111000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd375: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111110011000000000000000000110000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000000100000011100111110000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd376: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111111110000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111001111111111110000000000000000000001110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd377: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111111111111110000010111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000001111110000000001000000000000000011111111111110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd378: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111111111111111111111100011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110111010000000110000001110000000000000000010011110011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd379: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000001111111111111111111111111111111111011110101111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110000111111111000000000011000000000000000000110000111111111101111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd380: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000001111111111111111111111111111111111111000000001001111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000001110000011110000000000000000000001100011111111101110010110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd381: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000001111111111111111111111111111111111111000000011110000111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000001000000000000000000000000000000011100000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd382: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000011111111111111111111111111111111111101100011110011111111101111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000001010000000000000000000000000010011110000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd383: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111110011111101111111111110000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000011111110000000000111111110000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd384: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111110011110011111001111111111110111000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000011000000000000000000000000011101111111000000001110111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd385: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111000111111111001111111111111111100000000000000001111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101100000000000000100010000000000000000000001110101111110001000111110111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd386: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100000000000000111111111111111111111111111110001111111111111111111111111111111000000001000000000000001111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110011111111100000101011110111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd387: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010000000000000111111111111111111111111111110001111111111111111011111111111110000000010011100000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000100011111011001100010110010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd388: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110000000000000111111111111111111111111111100001111111111111111111111101000000000111100010000000000000000000000011111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000100000000000000000000000000000000001100000001100111111000000001111100001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd389: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000111111111111111111111111111100001111111111111111111111110011111011111111110000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000111100000111100100011110011001110000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd390: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000111111111110111111111111111100011111111111111111111111111111111100000011000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000010000000000000000000000010000000000000000000000000000000000000000001111001100000000011110000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd391: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000111111111111111111111111111100011111111111111111111111111111111111111111111111000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000010100000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd392: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000111111111111111111111111111000011111111111111111111111111111111111111111111111110000000001000000000000010000000000000001111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000001000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd393: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000011111111111111111111110000000011111111111111111111111111111111111111111111111111000000001100000000000000000000000000000000011111111111111111111100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000111100100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd394: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011000000000000011111111111111111111000000111111111111111111111111111111111111111111111111111111100000001110000000000000000000000000000000000000011111111111111111100000000000000000000001111110000000000000001100000000000000000000000000000000000000000000000000000111111100000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd395: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000000000000011111111111011111111000001111111111111111111111111111111111111111111111111111111100000000111100000000000000000000000000000000000000000111111111111111110000000000000000001111111011000010000000010000000000000000000000000000000000000000000000000001100111000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd396: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000011111111111111110000000011111111111111111111111111111111111111111111111111111111100000000011100000000000000000000000000000000000000000000001111111111111111100000000001111000011100000000000000000000000000000000000000000000000000000000000000000000011111111111000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd397: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000011111111111001000000001111111111111111111111111111111111111111111111111111111111110000000001110000000000000000000000000000000000000000000000000001111111111111111110000000000001000000000000001000000000000011100000000000000000000000000000000000000111111110011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd398: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000001111111100000000000011111111111111111111111111111111111111111111111111111111111100000000000111000000000000000000000000000000000000000000000000000000011111111111111111110000000001000000000000000000011010010000000000000000000000000010000000000001111111111101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd399: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000111111111000000000111111111111111111111111111111111111111111111111111111111111100000000001111100000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000010101100000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd400: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000011111111111000111111111111111111111111111111111111111111111111111111111111111100000000000101110000000000000000000000000000000000000000000000000000000000000011111111111111111111100000000000000000000111000000000000000000000000000000000000001111111100001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd401: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111100000011010100110000000000000000000000000000000000000000000000000000000000001111100111111111111111111111100000000000000000000000000000000000000000000000000100001111111111000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd402: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000001111111111111111111111111111111111111111111111111111111111111111111111100000001100000000000000000000000000000000000000000000000000000000000000000011111111111011111111111111111111111000000000000000000000000000000000000000000000000111111111111000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd403: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000011111111111111111111111111111111111111111111111111111111111111111100000000100000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111100000000000000000000000000000000000000001111110011011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd404: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000001111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000011111001111111111111111110000011111111111111111110000000000000000000000000000000000011111000001010111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd405: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000001111000001111111111111111100000000000111111111111111111110000000000000000000000000000111111000011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd406: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111100000000000000000010000000000000000000000000000000000000000000000000011111100111101111111111110000000000000000001111111111111111111100000000000000000000000000100000010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd407: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000001111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000111101111111111111111111111000000000000001111100000001111111111111111111100000000000000000111100000010100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd408: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000111111111111111111111111111111111111111111111001111111111100010000000000000000000000000000000000000000000000000000000000000110111111111011111111111110000000000000000001100000000000011111111111111111111110000001111111000000100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd409: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000001111111111111111111111111111111111111111111001111111111000000100000000000000000000000000000000000000000000000000000000001111111111111111111111111000100000000000000000000000000000000000111111111111111111111110011000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd410: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000011111111111111111111111111111111111111111011111111111000000000000000000000000000000000000000000000000000000000000000111111111111101111111111110010000000000000000000000000000000000000000000111111111111111111111000000001111011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd411: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000011111111111111111111111111111111111111111001111111110000000000000000000000000000000000000000000000000000000000000011111111111110111111111111000000000000000000000000000000000000000000000000000000011111111111111111111000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd412: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd413: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000100111111111111111111111111111111111111111111111000000001000000000000000000000000000000000000000000000000000000111111111110111111111111000000000000000000000000000000000000000000000000000000000011100101111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd414: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000011010111111111111111111111111111111111111111110000000001000000000000000000000000000000000000000000000000000000000111111001111111111110000000000000000000000000000000000000000000000000000000000001111111000000111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd415: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000011111101111111111111111111111111111111111111100000000001000000000000000000000000000000000000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000000000000000001111111000000000011111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd416: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000011111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000011111111111000001111111000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd417: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000011111110100011010001000011111000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd418: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000111111111110011100000000100111100000000000001111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd419: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000011111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000001111111111000000000000001000110000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd420: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000011111111111000111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000000001011110111100000000000000011011100000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd421: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000011111111100000000111111111111111110000000000000000000000000000000000000000011000001100000011000000000000111111111111000000000000000000000000000000000000000000000000000000000001111100111000000000000000001011000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd422: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000011111100000000000000000000000111110000000000000000000000000000000000000000000000011110000111000000000001111111111110000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000100000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd423: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000011110000000000000000000000000001111000000000000000000000000000000000000001100000101000011100000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd424: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000011110000000000000000000001111100000000000011000000000000000000000000000000110000100000100000000001011111111111110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd425: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000011111110000000000000000000011111100000000011111000000000000000000000000000000011000000000000000000100111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd426: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000011111110000000000000000000000001111110011111110000000000000000000000000000000011000000000000000000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd427: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000001111111000000000000000000110111111011111111110000000000000000000000000000000010000000000000000100111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd428: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000111111111000000000000000000011111111111111111110000000000000000000000000000000000000000000000001011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd429: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111100000000000000000011111111111111111100000000000000000000000000000000000000000000000000111111111111000010000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd430: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000111100001000000000000000000000011111111111111100000000000000000000000000000000000000000000000011111111111110000001100000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd431: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111111111111111111111110110000000000000000000000000001111100000000000000000000011111111111111100000000000000000000000000000000000000000000100111111111111100000100000010000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd432: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111110110000000000000000000000000000100100000000000000000001111111111111111000000000000000010000000000000000000000000000011111111111110000001100000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd433: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000100000000001000000000000000000000000000000011111111111111110000000000000000110000000000000000000000000000111111111111000000011100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd434: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111110100001110100110000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000001111111111110010101111100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd435: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111110001111100000001110000000000000001000000000000111111111111111100000000000000000000000000000000000000000100111111111111100000100000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd436: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111110000101101111111111000000000000000000000000000000011111111111100000000000000000000000000000000000000000000011111111111110000000100000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd437: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111011111111111110000000000000000000000000000000000011111111110000000000000000000000000000000000000011000000111111111111000000010101100000001100000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd438: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111000000000000000000000000000000000000011111111110000000000000000000000000000000000000000011111111111111110000001111111111000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd439: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111011101111111111000000000000000000000000000000000000000011111111100000000000000000000000010000000000000001000111111111111100000001101100110000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd440: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000010011111111111100000000000000000000000000000000000000000001111110000000000000000000000000000000000000000010011111111111110000000101111111000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd441: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000111111111111000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd442: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd443: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd444: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000;
			9'd445: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111000000000000000000000000000000000000000000000000000000000000;
			9'd446: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000;
			9'd447: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111110000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000;
			9'd448: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000010110000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000000;
			9'd449: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000;
			9'd450: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000000000000000000000;
			9'd451: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000;
			9'd452: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000010000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000;
			9'd453: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111000000000000000000;
			9'd454: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000;
			9'd455: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000;
			9'd456: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111;
			9'd457: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110011100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111;
			9'd458: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000011110000000000000000000000000000000000000000000000110000001000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111;
			9'd459: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101111111111000000000000000000000000000000000000000000000100001100000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100110001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111;
			9'd460: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000001111100000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd461: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111100011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd462: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000001000000000000000000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111011101111111100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd463: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101001111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd464: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd465: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100101111111111110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd466: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd467: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd468: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd469: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd470: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd471: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd472: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd473: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd474: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd475: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd476: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd477: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000100000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110011111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd478: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			9'd479: q <= 640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111110000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			default : q <= 640'd0;
		endcase	
	end
	assign out = q;
endmodule